`ifndef TR_FILE_LIST__SV 
`define TR_FILE_LIST__SV



`include "btslice.sv"

 `include "btslice_seq_sequence_library.sv"
`endif
