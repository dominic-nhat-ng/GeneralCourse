module testbench;
endmodule

