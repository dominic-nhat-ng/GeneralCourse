
`ifndef BTCOIN_MON_2COV_CONNECT
`define BTCOIN_MON_2COV_CONNECT
class btcoin_mon_2cov_connect extends uvm_component;
   btcoin_cov cov;
   uvm_analysis_export # (btcoin) an_exp;
   `uvm_component_utils(btcoin_mon_2cov_connect)
   function new(string name="", uvm_component parent=null);
   	super.new(name, parent);
   endfunction: new

   virtual function void write(btcoin tr);
      cov.tr = tr;
      -> cov.cov_event;
   endfunction:write 
endclass: btcoin_mon_2cov_connect

`endif // BTCOIN_MON_2COV_CONNECT
