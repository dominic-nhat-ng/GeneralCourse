VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

LAYER NWELL
  TYPE MASTERSLICE ;
END NWELL

LAYER PO
  TYPE MASTERSLICE ;
END PO

LAYER CO
  TYPE CUT ;
END CO

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.152 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M1

LAYER VIA1
  TYPE CUT ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.152 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M2

LAYER VIA2
  TYPE CUT ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M3

LAYER VIA3
  TYPE CUT ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M4

LAYER VIA4
  TYPE CUT ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M5

LAYER VIA5
  TYPE CUT ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M6

LAYER VIA6
  TYPE CUT ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M7

LAYER VIA7
  TYPE CUT ;
END VIA7

LAYER M8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M8

LAYER VIA8
  TYPE CUT ;
END VIA8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 2.432 ;
  WIDTH 0.16 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.16 WRONGDIRECTION ;" ;
END M9

LAYER VIARDL
  TYPE CUT ;
END VIARDL

LAYER MRDL
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 4.864 ;
  WIDTH 2 ;
  PROPERTY LEF58_WIDTH "WIDTH 2 WRONGDIRECTION ;" ;
END MRDL

LAYER DNW
  TYPE MASTERSLICE ;
END DNW

LAYER DIFF
  TYPE MASTERSLICE ;
END DIFF

LAYER PIMP
  TYPE MASTERSLICE ;
END PIMP

LAYER NIMP
  TYPE MASTERSLICE ;
END NIMP

LAYER DIFF_18
  TYPE MASTERSLICE ;
END DIFF_18

LAYER PAD
  TYPE MASTERSLICE ;
END PAD

LAYER ESD_25
  TYPE MASTERSLICE ;
END ESD_25

LAYER SBLK
  TYPE MASTERSLICE ;
END SBLK

LAYER HVTIMP
  TYPE MASTERSLICE ;
END HVTIMP

LAYER LVTIMP
  TYPE MASTERSLICE ;
END LVTIMP

LAYER M1PIN
  TYPE MASTERSLICE ;
END M1PIN

LAYER M2PIN
  TYPE MASTERSLICE ;
END M2PIN

LAYER M3PIN
  TYPE MASTERSLICE ;
END M3PIN

LAYER M4PIN
  TYPE MASTERSLICE ;
END M4PIN

LAYER M5PIN
  TYPE MASTERSLICE ;
END M5PIN

LAYER M6PIN
  TYPE MASTERSLICE ;
END M6PIN

LAYER M7PIN
  TYPE MASTERSLICE ;
END M7PIN

LAYER M8PIN
  TYPE MASTERSLICE ;
END M8PIN

LAYER M9PIN
  TYPE MASTERSLICE ;
END M9PIN

LAYER MRDL9PIN
  TYPE MASTERSLICE ;
END MRDL9PIN

LAYER HOTNWL
  TYPE MASTERSLICE ;
END HOTNWL

LAYER DIOD
  TYPE MASTERSLICE ;
END DIOD

LAYER BJTDMY
  TYPE MASTERSLICE ;
END BJTDMY

LAYER RNW
  TYPE MASTERSLICE ;
END RNW

LAYER RMARK
  TYPE MASTERSLICE ;
END RMARK

LAYER prBoundary
  TYPE MASTERSLICE ;
END prBoundary

LAYER LOGO
  TYPE MASTERSLICE ;
END LOGO

LAYER IP
  TYPE MASTERSLICE ;
END IP

LAYER RM1
  TYPE MASTERSLICE ;
END RM1

LAYER RM2
  TYPE MASTERSLICE ;
END RM2

LAYER RM3
  TYPE MASTERSLICE ;
END RM3

LAYER RM4
  TYPE MASTERSLICE ;
END RM4

LAYER RM5
  TYPE MASTERSLICE ;
END RM5

LAYER RM6
  TYPE MASTERSLICE ;
END RM6

LAYER RM7
  TYPE MASTERSLICE ;
END RM7

LAYER RM8
  TYPE MASTERSLICE ;
END RM8

LAYER RM9
  TYPE MASTERSLICE ;
END RM9

LAYER DM1EXCL
  TYPE MASTERSLICE ;
END DM1EXCL

LAYER DM2EXCL
  TYPE MASTERSLICE ;
END DM2EXCL

LAYER DM3EXCL
  TYPE MASTERSLICE ;
END DM3EXCL

LAYER DM4EXCL
  TYPE MASTERSLICE ;
END DM4EXCL

LAYER DM5EXCL
  TYPE MASTERSLICE ;
END DM5EXCL

LAYER DM6EXCL
  TYPE MASTERSLICE ;
END DM6EXCL

LAYER DM7EXCL
  TYPE MASTERSLICE ;
END DM7EXCL

LAYER DM8EXCL
  TYPE MASTERSLICE ;
END DM8EXCL

LAYER DM9EXCL
  TYPE MASTERSLICE ;
END DM9EXCL

LAYER DIFF_25
  TYPE MASTERSLICE ;
END DIFF_25

LAYER DIFF_FM
  TYPE MASTERSLICE ;
END DIFF_FM

LAYER PO_FM
  TYPE MASTERSLICE ;
END PO_FM

VIA VIA12SQ_C
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA12SQ_C

VIA VIA12BAR1_C
  LAYER M1 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA1 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA12BAR1_C

VIA VIA12BAR2_C
  LAYER M1 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M2 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA12BAR2_C

VIA VIA12LG_C
  LAYER M1 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA12LG_C

VIA VIA12SQ
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA12SQ

VIA VIA12BAR1
  LAYER M1 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA1 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M2 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA12BAR1

VIA VIA12BAR2
  LAYER M1 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA12BAR2

VIA VIA12LG
  LAYER M1 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA12LG

VIA VIA23SQ_C
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA23SQ_C

VIA VIA23BAR1_C
  LAYER M2 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA2 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA23BAR1_C

VIA VIA23BAR2_C
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M3 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA23BAR2_C

VIA VIA23LG_C
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA23LG_C

VIA VIA23SQ
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA23SQ

VIA VIA23BAR1
  LAYER M2 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA2 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M3 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA23BAR1

VIA VIA23BAR2
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA23BAR2

VIA VIA23LG
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA23LG

VIA VIA34SQ_C
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA34SQ_C

VIA VIA34BAR1_C
  LAYER M3 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA3 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA34BAR1_C

VIA VIA34BAR2_C
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M4 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA34BAR2_C

VIA VIA34LG_C
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA34LG_C

VIA VIA34SQ
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA34SQ

VIA VIA34BAR1
  LAYER M3 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA3 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M4 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA34BAR1

VIA VIA34BAR2
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA34BAR2

VIA VIA34LG
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA34LG

VIA VIA45SQ_C
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA45SQ_C

VIA VIA45BAR1_C
  LAYER M4 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA4 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA45BAR1_C

VIA VIA45BAR2_C
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M5 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA45BAR2_C

VIA VIA45LG_C
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA45LG_C

VIA VIA45SQ
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA45SQ

VIA VIA45BAR1
  LAYER M4 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA4 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M5 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA45BAR1

VIA VIA45BAR2
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA45BAR2

VIA VIA45LG
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA45LG

VIA VIA56SQ_C
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA56SQ_C

VIA VIA56BAR1_C
  LAYER M5 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA5 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA56BAR1_C

VIA VIA56BAR2_C
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M6 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA56BAR2_C

VIA VIA56LG_C
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA56LG_C

VIA VIA56SQ
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA56SQ

VIA VIA56BAR1
  LAYER M5 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA5 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M6 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA56BAR1

VIA VIA56BAR2
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA56BAR2

VIA VIA56LG
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA56LG

VIA VIA67SQ_C
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M7 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA67SQ_C

VIA VIA67BAR1_C
  LAYER M6 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA6 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA67BAR1_C

VIA VIA67BAR2_C
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M7 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA67BAR2_C

VIA VIA67LG_C
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA67LG_C

VIA VIA67SQ
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA67SQ

VIA VIA67BAR1
  LAYER M6 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA6 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M7 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA67BAR1

VIA VIA67BAR2
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA67BAR2

VIA VIA67LG
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA67LG

VIA VIA78SQ_C
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M8 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA78SQ_C

VIA VIA78BAR1_C
  LAYER M7 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA7 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M8 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA78BAR1_C

VIA VIA78BAR2_C
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M8 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA78BAR2_C

VIA VIA78LG_C
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M8 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA78LG_C

VIA VIA78SQ
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M8 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA78SQ

VIA VIA78BAR1
  LAYER M7 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA7 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M8 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA78BAR1

VIA VIA78BAR2
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M8 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA78BAR2

VIA VIA78LG
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M8 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA78LG

VIA VIA89_C
  LAYER M8 ;
    RECT -0.095 -0.08 0.095 0.08 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M9 ;
    RECT -0.08 -0.095 0.08 0.095 ;
END VIA89_C

VIA VIA89
  LAYER M8 ;
    RECT -0.095 -0.08 0.095 0.08 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M9 ;
    RECT -0.095 -0.08 0.095 0.08 ;
END VIA89

VIA VIA9RDL
  LAYER M9 ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER VIARDL ;
    RECT -1 -1 1 1 ;
  LAYER MRDL ;
    RECT -1.5 -1.5 1.5 1.5 ;
END VIA9RDL

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.152 BY 1.672 ;
END unit

MACRO bit_slice
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 200 BY 68 ;
  SYMMETRY X Y ;
  PIN hclk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 197.42 66.824 197.476 66.88 ;
        RECT 196.08 67.944 196.136 68 ;
    END
  END hclk
  PIN lclk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 197.724 66.824 197.78 66.88 ;
        RECT 196.384 67.944 196.44 68 ;
    END
  END lclk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.9 66.824 195.956 66.88 ;
        RECT 198.208 67.944 198.264 68 ;
    END
  END reset
  PIN sin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.572 66.824 26.628 66.88 ;
        RECT 2.01 67.944 2.066 68 ;
    END
  END sin
  PIN data_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.028 66.824 198.084 66.88 ;
        RECT 196.688 67.944 196.744 68 ;
    END
  END data_valid
  PIN memory_sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.412 66.824 128.468 66.88 ;
        RECT 184.348 67.944 184.404 68 ;
    END
  END memory_sleep
  PIN shut_down_signals[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.948 66.824 2.004 66.88 ;
        RECT 196.992 67.944 197.048 68 ;
    END
  END shut_down_signals[1]
  PIN shut_down_signals[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.644 66.824 1.7 66.88 ;
        RECT 197.296 67.944 197.352 68 ;
    END
  END shut_down_signals[0]
  PIN isolation_signals[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.34 66.824 1.396 66.88 ;
        RECT 2.19 67.944 2.246 68 ;
    END
  END isolation_signals[1]
  PIN isolation_signals[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.036 66.824 1.092 66.88 ;
        RECT 2.494 67.944 2.55 68 ;
    END
  END isolation_signals[0]
  PIN retention_signals[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.788 66.824 198.844 66.88 ;
        RECT 197.6 67.944 197.656 68 ;
    END
  END retention_signals[1]
  PIN retention_signals[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.092 66.824 199.148 66.88 ;
        RECT 197.904 67.944 197.96 68 ;
    END
  END retention_signals[0]
  PIN scan_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.332 66.824 198.388 66.88 ;
        RECT 171.58 67.944 171.636 68 ;
    END
  END scan_enable
  PIN sipo_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.676 66.824 106.732 66.88 ;
        RECT 3.102 67.944 3.158 68 ;
    END
  END sipo_scan_in
  PIN piso_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.796 66.824 39.852 66.88 ;
        RECT 2.01 67.944 2.066 68 ;
    END
  END piso_scan_in
  PIN hv_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.804 66.824 146.86 66.88 ;
        RECT 142.092 67.944 142.148 68 ;
    END
  END hv_scan_in
  PIN lv_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.052 66.824 120.108 66.88 ;
        RECT 79.924 67.944 79.98 68 ;
    END
  END lv_scan_in
  PIN sipo_scan_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.932 66.824 186.988 66.88 ;
        RECT 198.512 67.944 198.568 68 ;
    END
  END sipo_scan_out
  PIN piso_scan_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.268 66.824 26.324 66.88 ;
        RECT 198.804 67.944 198.86 68 ;
    END
  END piso_scan_out
  PIN hv_scan_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.596 66.824 195.652 66.88 ;
        RECT 12.892 67.944 12.948 68 ;
    END
  END hv_scan_out
  PIN lv_scan_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.798 67.944 2.854 68 ;
      LAYER M4 ;
        RECT 1.644 66.824 1.7 66.88 ;
    END
  END lv_scan_out
  PIN sout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.556 66.824 173.612 66.88 ;
        RECT 133.732 67.944 133.788 68 ;
    END
  END sout
  PIN memory_ack
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.18 66.824 160.236 66.88 ;
        RECT 187.236 67.944 187.292 68 ;
    END
  END memory_ack
  PIN PG_ack_signals[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.932 67.944 186.988 68 ;
      LAYER M4 ;
        RECT 3.772 66.824 3.828 66.88 ;
    END
  END PG_ack_signals[1]
  PIN PG_ack_signals[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.732 66.824 0.788 66.88 ;
        RECT 133.428 67.944 133.484 68 ;
    END
  END PG_ack_signals[0]
  PIN VDDH
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M8 ;
        RECT 28.5 0 31.5 3 ;
        RECT 92.5 0 95.5 3 ;
        RECT 158.5 0 161.5 3 ;
        RECT 28.5 63.88 31.5 66.88 ;
        RECT 92.5 63.88 95.5 66.88 ;
        RECT 158.5 63.88 161.5 66.88 ;
    END
  END VDDH
  PIN VDDL
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M8 ;
        RECT 38.5 0 41.5 3 ;
        RECT 102.5 0 105.5 3 ;
        RECT 168.5 0 171.5 3 ;
        RECT 38.5 63.88 41.5 66.88 ;
        RECT 102.5 63.88 105.5 66.88 ;
        RECT 168.5 63.88 171.5 66.88 ;
    END
  END VDDL
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M8 ;
        RECT 33.5 0 36.5 3 ;
        RECT 97.5 0 100.5 3 ;
        RECT 163.5 0 166.5 3 ;
        RECT 33.5 63.88 36.5 66.88 ;
        RECT 97.5 63.88 100.5 66.88 ;
        RECT 163.5 63.88 166.5 66.88 ;
    END
  END VSS
  PIN piso_sw_out
    DIRECTION OUTPUT ;
    USE POWER ;
  END piso_sw_out
  PIN sipo_sw_out
    DIRECTION OUTPUT ;
    USE POWER ;
  END sipo_sw_out
  OBS
    LAYER M2 ;
      RECT 172.336 67 172.856 67.3 ;
      RECT 185.104 67 186.232 67.3 ;
      RECT 80.68 64.3 105.976 67.3 ;
      RECT 129.168 64.3 132.728 67.3 ;
      RECT 134.488 64.3 141.392 67.3 ;
      RECT 142.848 64.3 146.104 67.3 ;
      RECT 160.936 64.3 170.88 67.3 ;
      RECT 174.312 64.3 183.648 67.3 ;
      RECT 187.992 64.3 194.896 67.3 ;
      RECT 3.858 64.3 12.192 67.3 ;
      RECT 13.648 64.3 25.568 67.3 ;
      RECT 40.552 64.3 79.224 67.3 ;
      RECT 40.552 64.3 79.224 67.3 ;
      RECT 80.68 64.3 105.976 67.3 ;
      RECT 77.68 64.244 80.68 67.244 ;
      RECT 0.7 0.7 199.3 66.124 ;
      RECT 107.432 64.3 119.352 67.3 ;
      RECT 120.808 64.3 127.712 67.3 ;
      RECT 147.56 64.3 159.48 67.3 ;
      RECT 129.168 64.3 132.728 67.3 ;
      RECT 134.488 64.3 141.392 67.3 ;
      RECT 142.848 64.3 146.104 67.3 ;
      RECT 131.488 64.244 134.488 67.244 ;
      RECT 139.848 64.244 142.848 67.244 ;
      RECT 160.936 64.3 170.88 67.3 ;
      RECT 169.856 64.244 172.856 67.244 ;
      RECT 174.312 64.3 183.648 67.3 ;
      RECT 183.232 64.244 186.232 67.244 ;
      RECT 187.992 64.3 194.896 67.3 ;
      RECT 187.688 64.244 190.688 67.244 ;
      RECT 27.328 64.3 39.096 67.3 ;
      RECT 3.858 64.3 12.192 67.3 ;
      RECT 13.648 64.3 25.568 67.3 ;
      RECT 2.704 64.244 5.704 67.244 ;
      RECT 10.648 64.244 13.648 67.244 ;
      POLYGON 143.822 67.999 143.822 67.869 143.82 67.869 143.82 67.3 146.104 67.3 146.104 66.124 147.56 66.124 147.56 67.3 152.73 67.3 152.73 67.391 152.79 67.391 152.79 67.3 156.836 67.3 156.836 67.585 156.834 67.585 156.834 67.695 156.894 67.695 156.894 67.585 156.892 67.585 156.892 67.3 159.48 67.3 159.48 66.124 160.936 66.124 160.936 67.3 170.88 67.3 170.88 67.244 172.336 67.244 172.336 67.3 172.856 67.3 172.856 66.124 174.312 66.124 174.312 67.3 180.852 67.3 180.852 67.565 180.85 67.565 180.85 67.695 180.91 67.695 180.91 67.565 180.908 67.565 180.908 67.3 183.648 67.3 183.648 67.244 184.348 67.244 184.348 67.261 184.346 67.261 184.346 67.391 184.406 67.391 184.406 67.261 184.404 67.261 184.404 67.244 185.104 67.244 185.104 67.3 185.562 67.3 185.562 67.391 185.622 67.391 185.622 67.3 186.232 67.3 186.232 66.124 187.688 66.124 187.688 67.244 187.992 67.244 187.992 67.3 188.298 67.3 188.298 67.391 188.358 67.391 188.358 67.3 194.896 67.3 194.896 66.124 196.48 66.124 196.48 66.48 196.592 66.48 196.592 66.124 196.656 66.124 196.656 67.244 196.72 67.244 196.72 66.124 198.484 66.124 198.484 66.369 198.482 66.369 198.482 66.479 198.542 66.479 198.542 66.369 198.54 66.369 198.54 66.124 199.3 66.124 199.3 0.7 196.412 0.7 196.412 0.683 196.414 0.683 196.414 0.553 196.354 0.553 196.354 0.683 196.356 0.683 196.356 0.7 154.156 0.7 154.156 0.379 154.158 0.379 154.158 0.249 154.098 0.249 154.098 0.379 154.1 0.379 154.1 0.7 146.1 0.7 146.1 0.511 146.102 0.511 146.102 0.401 146.042 0.401 146.042 0.511 146.044 0.511 146.044 0.7 136.524 0.7 136.524 0.227 136.526 0.227 136.526 0.097 136.466 0.097 136.466 0.227 136.468 0.227 136.468 0.7 135.46 0.7 135.46 0.531 135.462 0.531 135.462 0.401 135.402 0.401 135.402 0.531 135.404 0.531 135.404 0.7 131.66 0.7 131.66 0.683 131.662 0.683 131.662 0.553 131.602 0.553 131.602 0.683 131.604 0.683 131.604 0.7 126.036 0.7 126.036 0.379 126.038 0.379 126.038 0.249 125.978 0.249 125.978 0.379 125.98 0.379 125.98 0.7 109.772 0.7 109.772 0.531 109.774 0.531 109.774 0.401 109.714 0.401 109.714 0.531 109.716 0.531 109.716 0.7 103.996 0.7 103.996 0.486 104.023 0.486 104.023 0.426 103.913 0.426 103.913 0.486 103.94 0.486 103.94 0.7 103.54 0.7 103.54 0.531 103.542 0.531 103.542 0.401 103.482 0.401 103.482 0.531 103.484 0.531 103.484 0.7 78.308 0.7 78.308 0.182 78.335 0.182 78.335 0.122 78.225 0.122 78.225 0.182 78.252 0.182 78.252 0.7 76.484 0.7 76.484 0.227 76.486 0.227 76.486 0.097 76.426 0.097 76.426 0.227 76.428 0.227 76.428 0.7 72.836 0.7 72.836 0.683 72.838 0.683 72.838 0.553 72.778 0.553 72.778 0.683 72.78 0.683 72.78 0.7 0.7 0.7 0.7 66.124 2.704 66.124 2.704 67.244 3.858 67.244 3.858 67.3 6.964 67.3 6.964 67.565 6.962 67.565 6.962 67.695 7.022 67.695 7.022 67.565 7.02 67.565 7.02 67.3 12.192 67.3 12.192 67.244 13.648 67.244 13.648 67.3 25.568 67.3 25.568 66.124 27.328 66.124 27.328 67.3 29.762 67.3 29.762 67.391 29.822 67.391 29.822 67.3 39.096 67.3 39.096 66.124 40.552 66.124 40.552 67.3 79.012 67.3 79.012 67.565 79.01 67.565 79.01 67.695 79.07 67.695 79.07 67.565 79.068 67.565 79.068 67.3 79.224 67.3 79.224 67.244 80.68 67.244 80.68 67.3 105.976 67.3 105.976 66.124 106.98 66.124 106.98 66.197 106.978 66.197 106.978 66.327 107.038 66.327 107.038 66.197 107.036 66.197 107.036 66.124 107.432 66.124 107.432 67.3 119.352 67.3 119.352 66.124 120.808 66.124 120.808 67.3 127.712 67.3 127.712 66.124 129.168 66.124 129.168 67.3 130.996 67.3 130.996 67.869 130.994 67.869 130.994 67.999 131.054 67.999 131.054 67.869 131.052 67.869 131.052 67.3 132.728 67.3 132.728 67.244 134.488 67.244 134.488 67.3 137.074 67.3 137.074 67.391 137.134 67.391 137.134 67.3 141.392 67.3 141.392 67.244 142.848 67.244 142.848 67.3 143.764 67.3 143.764 67.869 143.762 67.869 143.762 67.999 ;
      POLYGON 127.862 67.999 127.862 67.889 127.86 67.889 127.86 67.58 127.804 67.58 127.804 67.889 127.802 67.889 127.802 67.999 ;
      POLYGON 120.718 67.999 120.718 67.869 120.716 67.869 120.716 66.479 120.718 66.479 120.718 66.369 120.658 66.369 120.658 66.479 120.66 66.479 120.66 67.869 120.658 67.869 120.658 67.999 ;
      POLYGON 198.694 67.695 198.694 67.585 198.692 67.585 198.692 66.347 198.694 66.347 198.694 66.217 198.634 66.217 198.634 66.347 198.636 66.347 198.636 67.585 198.634 67.585 198.634 67.695 ;
      RECT 120.354 67.124 120.414 67.391 ;
    LAYER M4 ;
      RECT 0.7 66.124 0.944 67.3 ;
      RECT 2.4 66.124 3.072 67.3 ;
      RECT 4.528 64.3 199.3 67.3 ;
      RECT 0.7 0.7 199.3 66.124 ;
      POLYGON 198.694 67.999 198.694 67.889 198.692 67.889 198.692 67.3 199.3 67.3 199.3 0.7 162.82 0.7 162.82 0.511 162.822 0.511 162.822 0.401 162.762 0.401 162.762 0.511 162.764 0.511 162.764 0.7 157.956 0.7 157.956 0.207 157.958 0.207 157.958 0.097 157.898 0.097 157.898 0.207 157.9 0.207 157.9 0.7 123.3 0.7 123.3 0.207 123.302 0.207 123.302 0.097 123.242 0.097 123.242 0.207 123.244 0.207 123.244 0.7 116.916 0.7 116.916 0.511 116.918 0.511 116.918 0.401 116.858 0.401 116.858 0.511 116.86 0.511 116.86 0.7 104.148 0.7 104.148 0.207 104.15 0.207 104.15 0.097 104.09 0.097 104.09 0.207 104.092 0.207 104.092 0.7 58.852 0.7 58.852 0.511 58.854 0.511 58.854 0.401 58.794 0.401 58.794 0.511 58.796 0.511 58.796 0.7 0.7 0.7 0.7 67.3 0.944 67.3 0.944 66.124 2.4 66.124 2.4 67.3 3.072 67.3 3.072 66.124 3.162 66.124 3.162 66.175 3.222 66.175 3.222 66.124 4.528 66.124 4.528 67.3 19.58 67.3 19.58 67.889 19.578 67.889 19.578 67.999 19.638 67.999 19.638 67.889 19.636 67.889 19.636 67.3 127.498 67.3 127.498 67.391 127.5 67.391 127.5 67.889 127.498 67.889 127.498 67.999 127.558 67.999 127.558 67.889 127.556 67.889 127.556 67.391 127.558 67.391 127.558 67.3 195.9 67.3 195.9 67.889 195.898 67.889 195.898 67.999 195.958 67.999 195.958 67.889 195.956 67.889 195.956 67.3 196.508 67.3 196.508 67.889 196.506 67.889 196.506 67.999 196.566 67.999 196.566 67.889 196.564 67.889 196.564 67.3 198.028 67.3 198.028 67.889 198.026 67.889 198.026 67.999 198.086 67.999 198.086 67.889 198.084 67.889 198.084 67.3 198.636 67.3 198.636 67.889 198.634 67.889 198.634 67.999 ;
      POLYGON 150.662 67.999 150.662 67.889 150.66 67.889 150.66 67.695 150.662 67.695 150.662 67.585 150.602 67.585 150.602 67.695 150.604 67.695 150.604 67.889 150.602 67.889 150.602 67.999 ;
      RECT 85.242 0.244 85.302 0.511 ;
    LAYER M8 ;
      RECT 32.2 63.18 32.8 67.3 ;
      RECT 37.2 63.18 37.8 67.3 ;
      RECT 96.2 63.18 96.8 67.3 ;
      RECT 101.2 63.18 101.8 67.3 ;
      RECT 162.2 63.18 162.8 67.3 ;
      RECT 167.2 63.18 167.8 67.3 ;
      RECT 32.2 0.7 32.8 3.7 ;
      RECT 37.2 0.7 37.8 3.7 ;
      RECT 96.2 0.7 96.8 3.7 ;
      RECT 101.2 0.7 101.8 3.7 ;
      RECT 162.2 0.7 162.8 3.7 ;
      RECT 167.2 0.7 167.8 3.7 ;
      RECT 0.7 63.18 27.8 67.3 ;
      RECT 42.2 63.18 91.8 67.3 ;
      RECT 106.2 63.18 157.8 67.3 ;
      RECT 172.2 63.18 199.3 67.3 ;
      RECT 0.7 3.7 199.3 63.18 ;
      RECT 0.7 0.7 27.8 3.7 ;
      RECT 42.2 0.7 91.8 3.7 ;
      RECT 106.2 0.7 157.8 3.7 ;
      RECT 172.2 0.7 199.3 3.7 ;
    LAYER NWELL ;
      RECT 0.23 0.23 199.77 67.77 ;
    LAYER PO ;
      RECT 0.122 0.122 199.878 67.878 ;
    LAYER M1 ;
      POLYGON 143.847 67.974 143.847 67.914 143.717 67.914 143.717 67.919 131.099 67.919 131.099 67.914 130.969 67.914 130.969 67.974 131.099 67.974 131.099 67.969 143.717 67.969 143.717 67.974 ;
      POLYGON 120.743 67.974 120.743 67.914 120.613 67.914 120.613 67.919 12.995 67.919 12.995 67.914 12.865 67.914 12.865 67.974 12.995 67.974 12.995 67.969 120.613 67.969 120.613 67.974 ;
      POLYGON 2.273 67.974 2.273 67.914 2.143 67.914 2.143 67.919 1.443 67.919 1.443 67.914 1.313 67.914 1.313 67.974 1.443 67.974 1.443 67.969 2.143 67.969 2.143 67.974 ;
      POLYGON 2.125 67.822 2.125 67.717 2.095 67.717 2.095 67.665 6.917 67.665 6.917 67.67 7.047 67.67 7.047 67.61 6.917 67.61 6.917 67.615 2.045 67.615 2.045 67.717 2.015 67.717 2.015 67.822 ;
      POLYGON 180.935 67.67 180.935 67.61 180.805 67.61 180.805 67.615 79.115 67.615 79.115 67.61 78.985 67.61 78.985 67.67 79.115 67.67 79.115 67.665 180.805 67.665 180.805 67.67 ;
      POLYGON 2.507 67.518 2.507 67.513 184.401 67.513 184.401 67.411 184.451 67.411 184.451 67.361 185.517 67.361 185.517 67.366 185.647 67.366 185.647 67.306 185.517 67.306 185.517 67.311 184.451 67.311 184.451 67.306 184.321 67.306 184.321 67.411 184.351 67.411 184.351 67.463 2.507 67.463 2.507 67.458 2.377 67.458 2.377 67.518 ;
      POLYGON 137.159 67.366 137.159 67.306 137.029 67.306 137.029 67.311 120.459 67.311 120.459 67.306 120.329 67.306 120.329 67.366 120.459 67.366 120.459 67.361 137.029 67.361 137.029 67.366 ;
      RECT 0.75 0.75 199.25 67.25 ;
      RECT 71.081 0.735 141.871 3.736 ;
      POLYGON 199.25 67.25 199.25 0.75 141.871 0.75 141.871 0.73 141.741 0.73 141.741 0.735 71.211 0.735 71.211 0.73 71.081 0.73 71.081 0.75 0.75 0.75 0.75 67.25 ;
      POLYGON 196.439 0.638 196.439 0.578 196.309 0.578 196.309 0.583 131.707 0.583 131.707 0.578 131.577 0.578 131.577 0.638 131.707 0.638 131.707 0.633 196.309 0.633 196.309 0.638 ;
      POLYGON 72.883 0.638 72.883 0.633 83.625 0.633 83.625 0.481 103.437 0.481 103.437 0.486 103.567 0.486 103.567 0.426 103.437 0.426 103.437 0.431 83.575 0.431 83.575 0.583 72.883 0.583 72.883 0.578 72.753 0.578 72.753 0.638 ;
      POLYGON 135.487 0.486 135.487 0.426 135.357 0.426 135.357 0.431 109.819 0.431 109.819 0.426 109.689 0.426 109.689 0.486 109.819 0.486 109.819 0.481 135.357 0.481 135.357 0.486 ;
      POLYGON 154.183 0.334 154.183 0.274 154.053 0.274 154.053 0.279 126.083 0.279 126.083 0.274 125.953 0.274 125.953 0.334 126.083 0.334 126.083 0.329 154.053 0.329 154.053 0.334 ;
      POLYGON 136.551 0.182 136.551 0.122 136.421 0.122 136.421 0.127 76.531 0.127 76.531 0.122 76.401 0.122 76.401 0.182 76.531 0.182 76.531 0.177 136.421 0.177 136.421 0.182 ;
    LAYER VIA1 ;
      RECT 143.767 67.919 143.817 67.969 ;
      RECT 130.999 67.919 131.049 67.969 ;
      RECT 120.663 67.919 120.713 67.969 ;
      RECT 12.895 67.919 12.945 67.969 ;
      RECT 2.193 67.919 2.243 67.969 ;
      RECT 1.343 67.919 1.393 67.969 ;
      RECT 2.045 67.767 2.095 67.817 ;
      RECT 180.855 67.615 180.905 67.665 ;
      RECT 79.015 67.615 79.065 67.665 ;
      RECT 6.967 67.615 7.017 67.665 ;
      RECT 2.407 67.463 2.457 67.513 ;
      RECT 185.567 67.311 185.617 67.361 ;
      RECT 184.351 67.311 184.401 67.361 ;
      RECT 137.079 67.311 137.129 67.361 ;
      RECT 120.359 67.311 120.409 67.361 ;
      RECT 2.013 67.159 2.063 67.209 ;
      RECT 198.791 67.007 198.841 67.057 ;
      RECT 197.575 67.007 197.625 67.057 ;
      RECT 186.935 67.007 186.985 67.057 ;
      RECT 196.967 66.551 197.017 66.601 ;
      RECT 2.559 66.551 2.609 66.601 ;
      RECT 1.039 66.551 1.089 66.601 ;
      RECT 198.639 66.247 198.689 66.297 ;
      RECT 106.983 66.247 107.033 66.297 ;
      RECT 39.799 66.095 39.849 66.145 ;
      RECT 141.791 0.735 141.841 0.785 ;
      RECT 71.111 0.735 71.161 0.785 ;
      RECT 196.359 0.583 196.409 0.633 ;
      RECT 131.607 0.583 131.657 0.633 ;
      RECT 72.783 0.583 72.833 0.633 ;
      RECT 135.407 0.431 135.457 0.481 ;
      RECT 109.719 0.431 109.769 0.481 ;
      RECT 103.487 0.431 103.537 0.481 ;
      RECT 154.103 0.279 154.153 0.329 ;
      RECT 125.983 0.279 126.033 0.329 ;
      RECT 136.471 0.127 136.521 0.177 ;
      RECT 76.431 0.127 76.481 0.177 ;
    LAYER VIA2 ;
      RECT 198.791 67.919 198.841 67.969 ;
      RECT 197.907 67.919 197.957 67.969 ;
      RECT 196.359 67.919 196.409 67.969 ;
      RECT 196.055 67.919 196.105 67.969 ;
      RECT 184.351 67.919 184.401 67.969 ;
      RECT 127.807 67.919 127.857 67.969 ;
      RECT 198.639 67.615 198.689 67.665 ;
      RECT 197.271 67.615 197.321 67.665 ;
      RECT 156.839 67.615 156.889 67.665 ;
      RECT 198.487 67.311 198.537 67.361 ;
      RECT 188.303 67.311 188.353 67.361 ;
      RECT 152.735 67.311 152.785 67.361 ;
      RECT 133.735 67.311 133.785 67.361 ;
      RECT 133.431 67.311 133.481 67.361 ;
      RECT 120.359 67.311 120.409 67.361 ;
      RECT 29.767 67.311 29.817 67.361 ;
      RECT 197.423 66.703 197.473 66.753 ;
      RECT 186.935 66.703 186.985 66.753 ;
      RECT 173.559 66.703 173.609 66.753 ;
      RECT 146.807 66.703 146.857 66.753 ;
      RECT 106.527 66.703 106.577 66.753 ;
      RECT 1.647 66.703 1.697 66.753 ;
      RECT 199.095 66.399 199.145 66.449 ;
      RECT 198.487 66.399 198.537 66.449 ;
      RECT 197.727 66.399 197.777 66.449 ;
      RECT 196.511 66.399 196.561 66.449 ;
      RECT 160.183 66.399 160.233 66.449 ;
      RECT 120.663 66.399 120.713 66.449 ;
      RECT 120.055 66.399 120.105 66.449 ;
      RECT 198.183 66.095 198.233 66.145 ;
      RECT 195.903 66.095 195.953 66.145 ;
      RECT 187.239 66.095 187.289 66.145 ;
      RECT 146.047 0.431 146.097 0.481 ;
      RECT 103.943 0.431 103.993 0.481 ;
      RECT 78.255 0.127 78.305 0.177 ;
    LAYER M3 ;
      RECT 198.604 67.914 198.871 67.974 ;
      RECT 197.844 67.914 198.111 67.974 ;
      RECT 196.324 67.914 196.591 67.974 ;
      RECT 195.868 67.914 196.135 67.974 ;
      POLYGON 184.431 67.974 184.431 67.914 184.321 67.914 184.321 67.916 127.887 67.916 127.887 67.914 127.777 67.914 127.777 67.974 127.887 67.974 127.887 67.972 184.321 67.972 184.321 67.974 ;
      POLYGON 127.583 67.974 127.583 67.914 127.473 67.914 127.473 67.916 19.663 67.916 19.663 67.914 19.553 67.914 19.553 67.974 19.663 67.974 19.663 67.972 127.473 67.972 127.473 67.974 ;
      POLYGON 198.719 67.67 198.719 67.61 198.609 67.61 198.609 67.612 197.351 67.612 197.351 67.61 197.241 67.61 197.241 67.67 197.351 67.67 197.351 67.668 198.609 67.668 198.609 67.67 ;
      POLYGON 156.919 67.67 156.919 67.61 156.809 67.61 156.809 67.612 150.687 67.612 150.687 67.61 150.577 67.61 150.577 67.67 150.687 67.67 150.687 67.668 156.809 67.668 156.809 67.67 ;
      POLYGON 198.567 67.366 198.567 67.306 198.457 67.306 198.457 67.308 188.383 67.308 188.383 67.306 188.273 67.306 188.273 67.366 188.383 67.366 188.383 67.364 198.457 67.364 198.457 67.366 ;
      POLYGON 152.815 67.366 152.815 67.306 152.705 67.306 152.705 67.308 133.815 67.308 133.815 67.306 133.705 67.306 133.705 67.366 133.815 67.366 133.815 67.364 152.705 67.364 152.705 67.366 ;
      POLYGON 133.511 67.366 133.511 67.306 133.401 67.306 133.401 67.308 127.583 67.308 127.583 67.306 127.473 67.306 127.473 67.366 127.583 67.366 127.583 67.364 133.401 67.364 133.401 67.366 ;
      POLYGON 120.439 67.366 120.439 67.306 120.329 67.306 120.329 67.308 29.847 67.308 29.847 67.306 29.737 67.306 29.737 67.366 29.847 67.366 29.847 67.364 120.329 67.364 120.329 67.366 ;
      RECT 0.7 0.7 199.3 67.3 ;
      POLYGON 199.3 67.3 199.3 0.7 145.492 0.7 145.492 0.484 146.017 0.484 146.017 0.486 146.127 0.486 146.127 0.426 146.017 0.426 146.017 0.428 145.436 0.428 145.436 0.7 0.7 0.7 0.7 67.3 ;
      POLYGON 103.998 0.511 103.998 0.401 103.938 0.401 103.938 0.428 85.327 0.428 85.327 0.426 85.217 0.426 85.217 0.486 85.327 0.486 85.327 0.484 103.938 0.484 103.938 0.511 ;
      POLYGON 78.31 0.207 78.31 0.18 104.065 0.18 104.065 0.182 104.175 0.182 104.175 0.122 104.065 0.122 104.065 0.124 78.31 0.124 78.31 0.097 78.25 0.097 78.25 0.207 ;
      POLYGON 157.983 0.182 157.983 0.122 157.873 0.122 157.873 0.124 123.327 0.124 123.327 0.122 123.217 0.122 123.217 0.182 123.327 0.182 123.327 0.18 157.873 0.18 157.873 0.182 ;
    LAYER VIA3 ;
      RECT 198.639 67.919 198.689 67.969 ;
      RECT 198.031 67.919 198.081 67.969 ;
      RECT 196.511 67.919 196.561 67.969 ;
      RECT 195.903 67.919 195.953 67.969 ;
      RECT 127.503 67.919 127.553 67.969 ;
      RECT 19.583 67.919 19.633 67.969 ;
      RECT 150.607 67.615 150.657 67.665 ;
      RECT 127.503 67.311 127.553 67.361 ;
      RECT 1.647 67.007 1.697 67.057 ;
      RECT 3.775 66.095 3.825 66.145 ;
      RECT 3.167 66.095 3.217 66.145 ;
      RECT 85.247 0.431 85.297 0.481 ;
      RECT 157.903 0.127 157.953 0.177 ;
      RECT 123.247 0.127 123.297 0.177 ;
      RECT 104.095 0.127 104.145 0.177 ;
    LAYER VIA4 ;
      RECT 150.607 67.919 150.657 67.969 ;
      RECT 3.167 66.095 3.217 66.145 ;
      RECT 162.767 0.431 162.817 0.481 ;
      RECT 116.863 0.431 116.913 0.481 ;
      RECT 85.247 0.431 85.297 0.481 ;
      RECT 58.799 0.431 58.849 0.481 ;
    LAYER M5 ;
      POLYGON 150.687 67.974 150.687 67.914 150.577 67.914 150.577 67.916 108.127 67.916 108.127 67.914 108.017 67.914 108.017 67.974 108.127 67.974 108.127 67.972 150.577 67.972 150.577 67.974 ;
      RECT 0.7 0.7 199.3 67.3 ;
      POLYGON 162.847 0.486 162.847 0.426 162.737 0.426 162.737 0.428 116.943 0.428 116.943 0.426 116.833 0.426 116.833 0.486 116.943 0.486 116.943 0.484 162.737 0.484 162.737 0.486 ;
      POLYGON 85.327 0.486 85.327 0.426 85.217 0.426 85.217 0.428 58.879 0.428 58.879 0.426 58.769 0.426 58.769 0.486 58.879 0.486 58.879 0.484 85.217 0.484 85.217 0.486 ;
    LAYER VIA5 ;
      RECT 108.047 67.919 108.097 67.969 ;
    LAYER M6 ;
      RECT 0.7 0.7 199.3 67.3 ;
      POLYGON 108.102 67.999 108.102 67.889 108.1 67.889 108.1 67.3 199.3 67.3 199.3 0.7 0.7 0.7 0.7 67.3 108.044 67.3 108.044 67.889 108.042 67.889 108.042 67.999 ;
    LAYER M7 ;
      RECT 0.7 0.7 199.3 67.3 ;
    LAYER VIA7 ;
      RECT 166.415 65.183 166.465 65.233 ;
      RECT 166.295 65.183 166.345 65.233 ;
      RECT 166.175 65.183 166.225 65.233 ;
      RECT 166.055 65.183 166.105 65.233 ;
      RECT 165.935 65.183 165.985 65.233 ;
      RECT 165.815 65.183 165.865 65.233 ;
      RECT 165.695 65.183 165.745 65.233 ;
      RECT 165.575 65.183 165.625 65.233 ;
      RECT 165.455 65.183 165.505 65.233 ;
      RECT 165.335 65.183 165.385 65.233 ;
      RECT 165.215 65.183 165.265 65.233 ;
      RECT 165.095 65.183 165.145 65.233 ;
      RECT 164.975 65.183 165.025 65.233 ;
      RECT 164.855 65.183 164.905 65.233 ;
      RECT 164.735 65.183 164.785 65.233 ;
      RECT 164.615 65.183 164.665 65.233 ;
      RECT 164.495 65.183 164.545 65.233 ;
      RECT 164.375 65.183 164.425 65.233 ;
      RECT 164.255 65.183 164.305 65.233 ;
      RECT 164.135 65.183 164.185 65.233 ;
      RECT 164.015 65.183 164.065 65.233 ;
      RECT 163.895 65.183 163.945 65.233 ;
      RECT 163.775 65.183 163.825 65.233 ;
      RECT 163.655 65.183 163.705 65.233 ;
      RECT 163.535 65.183 163.585 65.233 ;
      RECT 100.415 65.183 100.465 65.233 ;
      RECT 100.295 65.183 100.345 65.233 ;
      RECT 100.175 65.183 100.225 65.233 ;
      RECT 100.055 65.183 100.105 65.233 ;
      RECT 99.935 65.183 99.985 65.233 ;
      RECT 99.815 65.183 99.865 65.233 ;
      RECT 99.695 65.183 99.745 65.233 ;
      RECT 99.575 65.183 99.625 65.233 ;
      RECT 99.455 65.183 99.505 65.233 ;
      RECT 99.335 65.183 99.385 65.233 ;
      RECT 99.215 65.183 99.265 65.233 ;
      RECT 99.095 65.183 99.145 65.233 ;
      RECT 98.975 65.183 99.025 65.233 ;
      RECT 98.855 65.183 98.905 65.233 ;
      RECT 98.735 65.183 98.785 65.233 ;
      RECT 98.615 65.183 98.665 65.233 ;
      RECT 98.495 65.183 98.545 65.233 ;
      RECT 98.375 65.183 98.425 65.233 ;
      RECT 98.255 65.183 98.305 65.233 ;
      RECT 98.135 65.183 98.185 65.233 ;
      RECT 98.015 65.183 98.065 65.233 ;
      RECT 97.895 65.183 97.945 65.233 ;
      RECT 97.775 65.183 97.825 65.233 ;
      RECT 97.655 65.183 97.705 65.233 ;
      RECT 97.535 65.183 97.585 65.233 ;
      RECT 36.415 65.183 36.465 65.233 ;
      RECT 36.295 65.183 36.345 65.233 ;
      RECT 36.175 65.183 36.225 65.233 ;
      RECT 36.055 65.183 36.105 65.233 ;
      RECT 35.935 65.183 35.985 65.233 ;
      RECT 35.815 65.183 35.865 65.233 ;
      RECT 35.695 65.183 35.745 65.233 ;
      RECT 35.575 65.183 35.625 65.233 ;
      RECT 35.455 65.183 35.505 65.233 ;
      RECT 35.335 65.183 35.385 65.233 ;
      RECT 35.215 65.183 35.265 65.233 ;
      RECT 35.095 65.183 35.145 65.233 ;
      RECT 34.975 65.183 35.025 65.233 ;
      RECT 34.855 65.183 34.905 65.233 ;
      RECT 34.735 65.183 34.785 65.233 ;
      RECT 34.615 65.183 34.665 65.233 ;
      RECT 34.495 65.183 34.545 65.233 ;
      RECT 34.375 65.183 34.425 65.233 ;
      RECT 34.255 65.183 34.305 65.233 ;
      RECT 34.135 65.183 34.185 65.233 ;
      RECT 34.015 65.183 34.065 65.233 ;
      RECT 33.895 65.183 33.945 65.233 ;
      RECT 33.775 65.183 33.825 65.233 ;
      RECT 33.655 65.183 33.705 65.233 ;
      RECT 33.535 65.183 33.585 65.233 ;
      RECT 161.415 63.511 161.465 63.561 ;
      RECT 161.295 63.511 161.345 63.561 ;
      RECT 161.175 63.511 161.225 63.561 ;
      RECT 161.055 63.511 161.105 63.561 ;
      RECT 160.935 63.511 160.985 63.561 ;
      RECT 160.815 63.511 160.865 63.561 ;
      RECT 160.695 63.511 160.745 63.561 ;
      RECT 160.575 63.511 160.625 63.561 ;
      RECT 160.455 63.511 160.505 63.561 ;
      RECT 160.335 63.511 160.385 63.561 ;
      RECT 160.215 63.511 160.265 63.561 ;
      RECT 160.095 63.511 160.145 63.561 ;
      RECT 159.975 63.511 160.025 63.561 ;
      RECT 159.855 63.511 159.905 63.561 ;
      RECT 159.735 63.511 159.785 63.561 ;
      RECT 159.615 63.511 159.665 63.561 ;
      RECT 159.495 63.511 159.545 63.561 ;
      RECT 159.375 63.511 159.425 63.561 ;
      RECT 159.255 63.511 159.305 63.561 ;
      RECT 159.135 63.511 159.185 63.561 ;
      RECT 159.015 63.511 159.065 63.561 ;
      RECT 158.895 63.511 158.945 63.561 ;
      RECT 158.775 63.511 158.825 63.561 ;
      RECT 158.655 63.511 158.705 63.561 ;
      RECT 158.535 63.511 158.585 63.561 ;
      RECT 95.415 63.511 95.465 63.561 ;
      RECT 95.295 63.511 95.345 63.561 ;
      RECT 95.175 63.511 95.225 63.561 ;
      RECT 95.055 63.511 95.105 63.561 ;
      RECT 94.935 63.511 94.985 63.561 ;
      RECT 94.815 63.511 94.865 63.561 ;
      RECT 94.695 63.511 94.745 63.561 ;
      RECT 94.575 63.511 94.625 63.561 ;
      RECT 94.455 63.511 94.505 63.561 ;
      RECT 94.335 63.511 94.385 63.561 ;
      RECT 94.215 63.511 94.265 63.561 ;
      RECT 94.095 63.511 94.145 63.561 ;
      RECT 93.975 63.511 94.025 63.561 ;
      RECT 93.855 63.511 93.905 63.561 ;
      RECT 93.735 63.511 93.785 63.561 ;
      RECT 93.615 63.511 93.665 63.561 ;
      RECT 93.495 63.511 93.545 63.561 ;
      RECT 93.375 63.511 93.425 63.561 ;
      RECT 93.255 63.511 93.305 63.561 ;
      RECT 93.135 63.511 93.185 63.561 ;
      RECT 93.015 63.511 93.065 63.561 ;
      RECT 92.895 63.511 92.945 63.561 ;
      RECT 92.775 63.511 92.825 63.561 ;
      RECT 92.655 63.511 92.705 63.561 ;
      RECT 92.535 63.511 92.585 63.561 ;
      RECT 31.415 63.511 31.465 63.561 ;
      RECT 31.295 63.511 31.345 63.561 ;
      RECT 31.175 63.511 31.225 63.561 ;
      RECT 31.055 63.511 31.105 63.561 ;
      RECT 30.935 63.511 30.985 63.561 ;
      RECT 30.815 63.511 30.865 63.561 ;
      RECT 30.695 63.511 30.745 63.561 ;
      RECT 30.575 63.511 30.625 63.561 ;
      RECT 30.455 63.511 30.505 63.561 ;
      RECT 30.335 63.511 30.385 63.561 ;
      RECT 30.215 63.511 30.265 63.561 ;
      RECT 30.095 63.511 30.145 63.561 ;
      RECT 29.975 63.511 30.025 63.561 ;
      RECT 29.855 63.511 29.905 63.561 ;
      RECT 29.735 63.511 29.785 63.561 ;
      RECT 29.615 63.511 29.665 63.561 ;
      RECT 29.495 63.511 29.545 63.561 ;
      RECT 29.375 63.511 29.425 63.561 ;
      RECT 29.255 63.511 29.305 63.561 ;
      RECT 29.135 63.511 29.185 63.561 ;
      RECT 29.015 63.511 29.065 63.561 ;
      RECT 28.895 63.511 28.945 63.561 ;
      RECT 28.775 63.511 28.825 63.561 ;
      RECT 28.655 63.511 28.705 63.561 ;
      RECT 28.535 63.511 28.585 63.561 ;
      RECT 95.415 3.319 95.465 3.369 ;
      RECT 95.295 3.319 95.345 3.369 ;
      RECT 95.175 3.319 95.225 3.369 ;
      RECT 95.055 3.319 95.105 3.369 ;
      RECT 94.935 3.319 94.985 3.369 ;
      RECT 94.815 3.319 94.865 3.369 ;
      RECT 94.695 3.319 94.745 3.369 ;
      RECT 94.575 3.319 94.625 3.369 ;
      RECT 94.455 3.319 94.505 3.369 ;
      RECT 94.335 3.319 94.385 3.369 ;
      RECT 94.215 3.319 94.265 3.369 ;
      RECT 94.095 3.319 94.145 3.369 ;
      RECT 93.975 3.319 94.025 3.369 ;
      RECT 93.855 3.319 93.905 3.369 ;
      RECT 93.735 3.319 93.785 3.369 ;
      RECT 93.615 3.319 93.665 3.369 ;
      RECT 93.495 3.319 93.545 3.369 ;
      RECT 93.375 3.319 93.425 3.369 ;
      RECT 93.255 3.319 93.305 3.369 ;
      RECT 93.135 3.319 93.185 3.369 ;
      RECT 93.015 3.319 93.065 3.369 ;
      RECT 92.895 3.319 92.945 3.369 ;
      RECT 92.775 3.319 92.825 3.369 ;
      RECT 92.655 3.319 92.705 3.369 ;
      RECT 92.535 3.319 92.585 3.369 ;
      RECT 166.415 1.647 166.465 1.697 ;
      RECT 166.295 1.647 166.345 1.697 ;
      RECT 166.175 1.647 166.225 1.697 ;
      RECT 166.055 1.647 166.105 1.697 ;
      RECT 165.935 1.647 165.985 1.697 ;
      RECT 165.815 1.647 165.865 1.697 ;
      RECT 165.695 1.647 165.745 1.697 ;
      RECT 165.575 1.647 165.625 1.697 ;
      RECT 165.455 1.647 165.505 1.697 ;
      RECT 165.335 1.647 165.385 1.697 ;
      RECT 165.215 1.647 165.265 1.697 ;
      RECT 165.095 1.647 165.145 1.697 ;
      RECT 164.975 1.647 165.025 1.697 ;
      RECT 164.855 1.647 164.905 1.697 ;
      RECT 164.735 1.647 164.785 1.697 ;
      RECT 164.615 1.647 164.665 1.697 ;
      RECT 164.495 1.647 164.545 1.697 ;
      RECT 164.375 1.647 164.425 1.697 ;
      RECT 164.255 1.647 164.305 1.697 ;
      RECT 164.135 1.647 164.185 1.697 ;
      RECT 164.015 1.647 164.065 1.697 ;
      RECT 163.895 1.647 163.945 1.697 ;
      RECT 163.775 1.647 163.825 1.697 ;
      RECT 163.655 1.647 163.705 1.697 ;
      RECT 163.535 1.647 163.585 1.697 ;
      RECT 100.415 1.647 100.465 1.697 ;
      RECT 100.295 1.647 100.345 1.697 ;
      RECT 100.175 1.647 100.225 1.697 ;
      RECT 100.055 1.647 100.105 1.697 ;
      RECT 99.935 1.647 99.985 1.697 ;
      RECT 99.815 1.647 99.865 1.697 ;
      RECT 99.695 1.647 99.745 1.697 ;
      RECT 99.575 1.647 99.625 1.697 ;
      RECT 99.455 1.647 99.505 1.697 ;
      RECT 99.335 1.647 99.385 1.697 ;
      RECT 99.215 1.647 99.265 1.697 ;
      RECT 99.095 1.647 99.145 1.697 ;
      RECT 98.975 1.647 99.025 1.697 ;
      RECT 98.855 1.647 98.905 1.697 ;
      RECT 98.735 1.647 98.785 1.697 ;
      RECT 98.615 1.647 98.665 1.697 ;
      RECT 98.495 1.647 98.545 1.697 ;
      RECT 98.375 1.647 98.425 1.697 ;
      RECT 98.255 1.647 98.305 1.697 ;
      RECT 98.135 1.647 98.185 1.697 ;
      RECT 98.015 1.647 98.065 1.697 ;
      RECT 97.895 1.647 97.945 1.697 ;
      RECT 97.775 1.647 97.825 1.697 ;
      RECT 97.655 1.647 97.705 1.697 ;
      RECT 97.535 1.647 97.585 1.697 ;
      RECT 36.415 1.647 36.465 1.697 ;
      RECT 36.295 1.647 36.345 1.697 ;
      RECT 36.175 1.647 36.225 1.697 ;
      RECT 36.055 1.647 36.105 1.697 ;
      RECT 35.935 1.647 35.985 1.697 ;
      RECT 35.815 1.647 35.865 1.697 ;
      RECT 35.695 1.647 35.745 1.697 ;
      RECT 35.575 1.647 35.625 1.697 ;
      RECT 35.455 1.647 35.505 1.697 ;
      RECT 35.335 1.647 35.385 1.697 ;
      RECT 35.215 1.647 35.265 1.697 ;
      RECT 35.095 1.647 35.145 1.697 ;
      RECT 34.975 1.647 35.025 1.697 ;
      RECT 34.855 1.647 34.905 1.697 ;
      RECT 34.735 1.647 34.785 1.697 ;
      RECT 34.615 1.647 34.665 1.697 ;
      RECT 34.495 1.647 34.545 1.697 ;
      RECT 34.375 1.647 34.425 1.697 ;
      RECT 34.255 1.647 34.305 1.697 ;
      RECT 34.135 1.647 34.185 1.697 ;
      RECT 34.015 1.647 34.065 1.697 ;
      RECT 33.895 1.647 33.945 1.697 ;
      RECT 33.775 1.647 33.825 1.697 ;
      RECT 33.655 1.647 33.705 1.697 ;
      RECT 33.535 1.647 33.585 1.697 ;
    LAYER M9 ;
      RECT 0.5 0.5 199.5 67.5 ;
    LAYER MRDL ;
      RECT 2 2 198 66 ;
  END
END bit_slice

END LIBRARY
