`timescale 1ns/1ps;

`include "uvm_macros.svh"

import uvm_pkg::*;

module testbench;


endmodule
