class base_test extends uvm_test;

endclass
