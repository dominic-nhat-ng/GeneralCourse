VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

LAYER NWELL
  TYPE MASTERSLICE ;
END NWELL

LAYER PO
  TYPE MASTERSLICE ;
END PO

LAYER CO
  TYPE CUT ;
END CO

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.152 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M1

LAYER VIA1
  TYPE CUT ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.152 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M2

LAYER VIA2
  TYPE CUT ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M3

LAYER VIA3
  TYPE CUT ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M4

LAYER VIA4
  TYPE CUT ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M5

LAYER VIA5
  TYPE CUT ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M6

LAYER VIA6
  TYPE CUT ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M7

LAYER VIA7
  TYPE CUT ;
END VIA7

LAYER M8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M8

LAYER VIA8
  TYPE CUT ;
END VIA8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 2.432 ;
  WIDTH 0.16 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.16 WRONGDIRECTION ;" ;
END M9

LAYER VIARDL
  TYPE CUT ;
END VIARDL

LAYER MRDL
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 4.864 ;
  WIDTH 2 ;
  PROPERTY LEF58_WIDTH "WIDTH 2 WRONGDIRECTION ;" ;
END MRDL

LAYER DNW
  TYPE MASTERSLICE ;
END DNW

LAYER DIFF
  TYPE MASTERSLICE ;
END DIFF

LAYER PIMP
  TYPE MASTERSLICE ;
END PIMP

LAYER NIMP
  TYPE MASTERSLICE ;
END NIMP

LAYER DIFF_18
  TYPE MASTERSLICE ;
END DIFF_18

LAYER PAD
  TYPE MASTERSLICE ;
END PAD

LAYER ESD_25
  TYPE MASTERSLICE ;
END ESD_25

LAYER SBLK
  TYPE MASTERSLICE ;
END SBLK

LAYER HVTIMP
  TYPE MASTERSLICE ;
END HVTIMP

LAYER LVTIMP
  TYPE MASTERSLICE ;
END LVTIMP

LAYER M1PIN
  TYPE MASTERSLICE ;
END M1PIN

LAYER M2PIN
  TYPE MASTERSLICE ;
END M2PIN

LAYER M3PIN
  TYPE MASTERSLICE ;
END M3PIN

LAYER M4PIN
  TYPE MASTERSLICE ;
END M4PIN

LAYER M5PIN
  TYPE MASTERSLICE ;
END M5PIN

LAYER M6PIN
  TYPE MASTERSLICE ;
END M6PIN

LAYER M7PIN
  TYPE MASTERSLICE ;
END M7PIN

LAYER M8PIN
  TYPE MASTERSLICE ;
END M8PIN

LAYER M9PIN
  TYPE MASTERSLICE ;
END M9PIN

LAYER MRDL9PIN
  TYPE MASTERSLICE ;
END MRDL9PIN

LAYER HOTNWL
  TYPE MASTERSLICE ;
END HOTNWL

LAYER DIOD
  TYPE MASTERSLICE ;
END DIOD

LAYER BJTDMY
  TYPE MASTERSLICE ;
END BJTDMY

LAYER RNW
  TYPE MASTERSLICE ;
END RNW

LAYER RMARK
  TYPE MASTERSLICE ;
END RMARK

LAYER prBoundary
  TYPE MASTERSLICE ;
END prBoundary

LAYER LOGO
  TYPE MASTERSLICE ;
END LOGO

LAYER IP
  TYPE MASTERSLICE ;
END IP

LAYER RM1
  TYPE MASTERSLICE ;
END RM1

LAYER RM2
  TYPE MASTERSLICE ;
END RM2

LAYER RM3
  TYPE MASTERSLICE ;
END RM3

LAYER RM4
  TYPE MASTERSLICE ;
END RM4

LAYER RM5
  TYPE MASTERSLICE ;
END RM5

LAYER RM6
  TYPE MASTERSLICE ;
END RM6

LAYER RM7
  TYPE MASTERSLICE ;
END RM7

LAYER RM8
  TYPE MASTERSLICE ;
END RM8

LAYER RM9
  TYPE MASTERSLICE ;
END RM9

LAYER DM1EXCL
  TYPE MASTERSLICE ;
END DM1EXCL

LAYER DM2EXCL
  TYPE MASTERSLICE ;
END DM2EXCL

LAYER DM3EXCL
  TYPE MASTERSLICE ;
END DM3EXCL

LAYER DM4EXCL
  TYPE MASTERSLICE ;
END DM4EXCL

LAYER DM5EXCL
  TYPE MASTERSLICE ;
END DM5EXCL

LAYER DM6EXCL
  TYPE MASTERSLICE ;
END DM6EXCL

LAYER DM7EXCL
  TYPE MASTERSLICE ;
END DM7EXCL

LAYER DM8EXCL
  TYPE MASTERSLICE ;
END DM8EXCL

LAYER DM9EXCL
  TYPE MASTERSLICE ;
END DM9EXCL

LAYER DIFF_25
  TYPE MASTERSLICE ;
END DIFF_25

LAYER DIFF_FM
  TYPE MASTERSLICE ;
END DIFF_FM

LAYER PO_FM
  TYPE MASTERSLICE ;
END PO_FM

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA VIA12SQ_C
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA12SQ_C

VIA VIA12BAR1_C
  LAYER M1 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA1 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA12BAR1_C

VIA VIA12BAR2_C
  LAYER M1 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M2 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA12BAR2_C

VIA VIA12LG_C
  LAYER M1 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA12LG_C

VIA VIA12SQ
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA12SQ

VIA VIA12BAR1
  LAYER M1 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA1 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M2 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA12BAR1

VIA VIA12BAR2
  LAYER M1 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA12BAR2

VIA VIA12LG
  LAYER M1 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA12LG

VIA VIA23SQ_C
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA23SQ_C

VIA VIA23BAR1_C
  LAYER M2 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA2 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA23BAR1_C

VIA VIA23BAR2_C
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M3 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA23BAR2_C

VIA VIA23LG_C
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA23LG_C

VIA VIA23SQ
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA23SQ

VIA VIA23BAR1
  LAYER M2 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA2 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M3 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA23BAR1

VIA VIA23BAR2
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA23BAR2

VIA VIA23LG
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA23LG

VIA VIA34SQ_C
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA34SQ_C

VIA VIA34BAR1_C
  LAYER M3 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA3 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA34BAR1_C

VIA VIA34BAR2_C
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M4 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA34BAR2_C

VIA VIA34LG_C
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA34LG_C

VIA VIA34SQ
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA34SQ

VIA VIA34BAR1
  LAYER M3 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA3 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M4 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA34BAR1

VIA VIA34BAR2
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA34BAR2

VIA VIA34LG
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA34LG

VIA VIA45SQ_C
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA45SQ_C

VIA VIA45BAR1_C
  LAYER M4 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA4 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA45BAR1_C

VIA VIA45BAR2_C
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M5 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA45BAR2_C

VIA VIA45LG_C
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA45LG_C

VIA VIA45SQ
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA45SQ

VIA VIA45BAR1
  LAYER M4 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA4 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M5 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA45BAR1

VIA VIA45BAR2
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA45BAR2

VIA VIA45LG
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA45LG

VIA VIA56SQ_C
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA56SQ_C

VIA VIA56BAR1_C
  LAYER M5 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA5 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA56BAR1_C

VIA VIA56BAR2_C
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M6 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA56BAR2_C

VIA VIA56LG_C
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA56LG_C

VIA VIA56SQ
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA56SQ

VIA VIA56BAR1
  LAYER M5 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA5 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M6 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA56BAR1

VIA VIA56BAR2
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA56BAR2

VIA VIA56LG
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA56LG

VIA VIA67SQ_C
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M7 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA67SQ_C

VIA VIA67BAR1_C
  LAYER M6 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA6 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA67BAR1_C

VIA VIA67BAR2_C
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M7 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA67BAR2_C

VIA VIA67LG_C
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA67LG_C

VIA VIA67SQ
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA67SQ

VIA VIA67BAR1
  LAYER M6 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA6 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M7 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA67BAR1

VIA VIA67BAR2
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA67BAR2

VIA VIA67LG
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA67LG

VIA VIA78SQ_C
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M8 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA78SQ_C

VIA VIA78BAR1_C
  LAYER M7 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA7 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M8 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA78BAR1_C

VIA VIA78BAR2_C
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M8 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA78BAR2_C

VIA VIA78LG_C
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M8 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA78LG_C

VIA VIA78SQ
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M8 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA78SQ

VIA VIA78BAR1
  LAYER M7 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER VIA7 ;
    RECT -0.05 -0.025 0.05 0.025 ;
  LAYER M8 ;
    RECT -0.08 -0.03 0.08 0.03 ;
END VIA78BAR1

VIA VIA78BAR2
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M8 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA78BAR2

VIA VIA78LG
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M8 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA78LG

VIA VIA89_C
  LAYER M8 ;
    RECT -0.095 -0.08 0.095 0.08 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M9 ;
    RECT -0.08 -0.095 0.08 0.095 ;
END VIA89_C

VIA VIA89
  LAYER M8 ;
    RECT -0.095 -0.08 0.095 0.08 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M9 ;
    RECT -0.095 -0.08 0.095 0.08 ;
END VIA89

VIA VIA9RDL
  LAYER M9 ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER VIARDL ;
    RECT -1 -1 1 1 ;
  LAYER MRDL ;
    RECT -1.5 -1.5 1.5 1.5 ;
END VIA9RDL

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.152 BY 1.672 ;
END unit

MACRO bit_top
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 1638.912 BY 468.816 ;
  SYMMETRY X Y ;
  PIN hclk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 807.876 468.76 807.932 468.816 ;
    END
  END hclk
  PIN lclk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 810.916 468.76 810.972 468.816 ;
    END
  END lclk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 811.524 468.76 811.58 468.816 ;
    END
  END reset
  PIN data_in_serial
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 508.588 468.76 508.644 468.816 ;
    END
  END data_in_serial
  PIN data_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 807.572 468.76 807.628 468.816 ;
    END
  END data_valid
  PIN memory_sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 802.86 468.76 802.916 468.816 ;
    END
  END memory_sleep
  PIN shut_down_signals[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 613.62 468.76 613.676 468.816 ;
    END
  END shut_down_signals[1]
  PIN shut_down_signals[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1005.628 468.76 1005.684 468.816 ;
    END
  END shut_down_signals[0]
  PIN isolation_signals[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 808.484 468.76 808.54 468.816 ;
    END
  END isolation_signals[1]
  PIN isolation_signals[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 808.18 468.76 808.236 468.816 ;
    END
  END isolation_signals[0]
  PIN retention_signals[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 811.22 468.76 811.276 468.816 ;
    END
  END retention_signals[1]
  PIN retention_signals[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 810.612 468.76 810.668 468.816 ;
    END
  END retention_signals[0]
  PIN scan_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 776.108 468.76 776.164 468.816 ;
    END
  END scan_enable
  PIN sipo_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 722.604 468.76 722.66 468.816 ;
    END
  END sipo_scan_in
  PIN piso_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 923.244 468.76 923.3 468.816 ;
    END
  END piso_scan_in
  PIN hv_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.324 468.76 321.38 468.816 ;
    END
  END hv_scan_in
  PIN lv_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 695.852 468.76 695.908 468.816 ;
    END
  END lv_scan_in
  PIN sipo_scan_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 898.468 468.76 898.524 468.816 ;
    END
  END sipo_scan_out
  PIN piso_scan_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 785.684 468.76 785.74 468.816 ;
    END
  END piso_scan_out
  PIN hv_scan_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 650.556 468.76 650.612 468.816 ;
    END
  END hv_scan_out
  PIN lv_scan_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.548 468.76 11.604 468.816 ;
    END
  END lv_scan_out
  PIN sout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 611.036 468.76 611.092 468.816 ;
    END
  END sout[1]
  PIN sout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 544.916 468.76 544.972 468.816 ;
    END
  END sout[0]
  PIN memory_address[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.508 468.76 350.564 468.816 ;
    END
  END memory_address[3]
  PIN memory_address[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.332 468.76 219.388 468.816 ;
    END
  END memory_address[2]
  PIN memory_address[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 534.124 468.76 534.18 468.816 ;
    END
  END memory_address[1]
  PIN memory_address[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1197.908 468.76 1197.964 468.816 ;
    END
  END memory_address[0]
  PIN memory_ack
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1487.62 468.76 1487.676 468.816 ;
    END
  END memory_ack
  PIN PG_ack_signals[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.516 468.76 77.572 468.816 ;
    END
  END PG_ack_signals[3]
  PIN PG_ack_signals[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.444 468.76 26.5 468.816 ;
    END
  END PG_ack_signals[2]
  PIN PG_ack_signals[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1438.22 468.76 1438.276 468.816 ;
    END
  END PG_ack_signals[1]
  PIN PG_ack_signals[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1302.18 468.76 1302.236 468.816 ;
    END
  END PG_ack_signals[0]
  PIN VDDH
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M8 ;
        RECT 38.5 0 41.5 3 ;
        RECT 102.5 0 105.5 3 ;
        RECT 168.5 0 171.5 3 ;
        RECT 238.5 0 241.5 3 ;
        RECT 302.5 0 305.5 3 ;
        RECT 368.5 0 371.5 3 ;
        RECT 438.5 0 441.5 3 ;
        RECT 502.5 0 505.5 3 ;
        RECT 568.5 0 571.5 3 ;
        RECT 638.5 0 641.5 3 ;
        RECT 702.5 0 705.5 3 ;
        RECT 768.5 0 771.5 3 ;
        RECT 838.5 0 841.5 3 ;
        RECT 902.5 0 905.5 3 ;
        RECT 968.5 0 971.5 3 ;
        RECT 1038.5 0 1041.5 3 ;
        RECT 1102.5 0 1105.5 3 ;
        RECT 1168.5 0 1171.5 3 ;
        RECT 1238.5 0 1241.5 3 ;
        RECT 1302.5 0 1305.5 3 ;
        RECT 1368.5 0 1371.5 3 ;
        RECT 1438.5 0 1441.5 3 ;
        RECT 1502.5 0 1505.5 3 ;
        RECT 1568.5 0 1571.5 3 ;
        RECT 38.5 465.816 41.5 468.816 ;
        RECT 102.5 465.816 105.5 468.816 ;
        RECT 168.5 465.816 171.5 468.816 ;
        RECT 238.5 465.816 241.5 468.816 ;
        RECT 302.5 465.816 305.5 468.816 ;
        RECT 368.5 465.816 371.5 468.816 ;
        RECT 438.5 465.816 441.5 468.816 ;
        RECT 502.5 465.816 505.5 468.816 ;
        RECT 568.5 465.816 571.5 468.816 ;
        RECT 638.5 465.816 641.5 468.816 ;
        RECT 702.5 465.816 705.5 468.816 ;
        RECT 768.5 465.816 771.5 468.816 ;
        RECT 838.5 465.816 841.5 468.816 ;
        RECT 902.5 465.816 905.5 468.816 ;
        RECT 968.5 465.816 971.5 468.816 ;
        RECT 1038.5 465.816 1041.5 468.816 ;
        RECT 1102.5 465.816 1105.5 468.816 ;
        RECT 1168.5 465.816 1171.5 468.816 ;
        RECT 1238.5 465.816 1241.5 468.816 ;
        RECT 1302.5 465.816 1305.5 468.816 ;
        RECT 1368.5 465.816 1371.5 468.816 ;
        RECT 1438.5 465.816 1441.5 468.816 ;
        RECT 1502.5 465.816 1505.5 468.816 ;
        RECT 1568.5 465.816 1571.5 468.816 ;
    END
  END VDDH
  PIN VDDL
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M8 ;
        RECT 48.5 0 51.5 3 ;
        RECT 112.5 0 115.5 3 ;
        RECT 178.5 0 181.5 3 ;
        RECT 248.5 0 251.5 3 ;
        RECT 312.5 0 315.5 3 ;
        RECT 378.5 0 381.5 3 ;
        RECT 448.5 0 451.5 3 ;
        RECT 512.5 0 515.5 3 ;
        RECT 578.5 0 581.5 3 ;
        RECT 648.5 0 651.5 3 ;
        RECT 712.5 0 715.5 3 ;
        RECT 778.5 0 781.5 3 ;
        RECT 848.5 0 851.5 3 ;
        RECT 912.5 0 915.5 3 ;
        RECT 978.5 0 981.5 3 ;
        RECT 1048.5 0 1051.5 3 ;
        RECT 1112.5 0 1115.5 3 ;
        RECT 1178.5 0 1181.5 3 ;
        RECT 1248.5 0 1251.5 3 ;
        RECT 1312.5 0 1315.5 3 ;
        RECT 1378.5 0 1381.5 3 ;
        RECT 1448.5 0 1451.5 3 ;
        RECT 1512.5 0 1515.5 3 ;
        RECT 1578.5 0 1581.5 3 ;
        RECT 48.5 465.816 51.5 468.816 ;
        RECT 112.5 465.816 115.5 468.816 ;
        RECT 178.5 465.816 181.5 468.816 ;
        RECT 248.5 465.816 251.5 468.816 ;
        RECT 312.5 465.816 315.5 468.816 ;
        RECT 378.5 465.816 381.5 468.816 ;
        RECT 448.5 465.816 451.5 468.816 ;
        RECT 512.5 465.816 515.5 468.816 ;
        RECT 578.5 465.816 581.5 468.816 ;
        RECT 648.5 465.816 651.5 468.816 ;
        RECT 712.5 465.816 715.5 468.816 ;
        RECT 778.5 465.816 781.5 468.816 ;
        RECT 848.5 465.816 851.5 468.816 ;
        RECT 912.5 465.816 915.5 468.816 ;
        RECT 978.5 465.816 981.5 468.816 ;
        RECT 1048.5 465.816 1051.5 468.816 ;
        RECT 1112.5 465.816 1115.5 468.816 ;
        RECT 1178.5 465.816 1181.5 468.816 ;
        RECT 1248.5 465.816 1251.5 468.816 ;
        RECT 1312.5 465.816 1315.5 468.816 ;
        RECT 1378.5 465.816 1381.5 468.816 ;
        RECT 1448.5 465.816 1451.5 468.816 ;
        RECT 1512.5 465.816 1515.5 468.816 ;
        RECT 1578.5 465.816 1581.5 468.816 ;
    END
  END VDDL
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M8 ;
        RECT 43.5 0 46.5 3 ;
        RECT 107.5 0 110.5 3 ;
        RECT 173.5 0 176.5 3 ;
        RECT 243.5 0 246.5 3 ;
        RECT 307.5 0 310.5 3 ;
        RECT 373.5 0 376.5 3 ;
        RECT 443.5 0 446.5 3 ;
        RECT 507.5 0 510.5 3 ;
        RECT 573.5 0 576.5 3 ;
        RECT 643.5 0 646.5 3 ;
        RECT 707.5 0 710.5 3 ;
        RECT 773.5 0 776.5 3 ;
        RECT 843.5 0 846.5 3 ;
        RECT 907.5 0 910.5 3 ;
        RECT 973.5 0 976.5 3 ;
        RECT 1043.5 0 1046.5 3 ;
        RECT 1107.5 0 1110.5 3 ;
        RECT 1173.5 0 1176.5 3 ;
        RECT 1243.5 0 1246.5 3 ;
        RECT 1307.5 0 1310.5 3 ;
        RECT 1373.5 0 1376.5 3 ;
        RECT 1443.5 0 1446.5 3 ;
        RECT 1507.5 0 1510.5 3 ;
        RECT 1573.5 0 1576.5 3 ;
        RECT 43.5 465.816 46.5 468.816 ;
        RECT 107.5 465.816 110.5 468.816 ;
        RECT 173.5 465.816 176.5 468.816 ;
        RECT 243.5 465.816 246.5 468.816 ;
        RECT 307.5 465.816 310.5 468.816 ;
        RECT 373.5 465.816 376.5 468.816 ;
        RECT 443.5 465.816 446.5 468.816 ;
        RECT 507.5 465.816 510.5 468.816 ;
        RECT 573.5 465.816 576.5 468.816 ;
        RECT 643.5 465.816 646.5 468.816 ;
        RECT 707.5 465.816 710.5 468.816 ;
        RECT 773.5 465.816 776.5 468.816 ;
        RECT 843.5 465.816 846.5 468.816 ;
        RECT 907.5 465.816 910.5 468.816 ;
        RECT 973.5 465.816 976.5 468.816 ;
        RECT 1043.5 465.816 1046.5 468.816 ;
        RECT 1107.5 465.816 1110.5 468.816 ;
        RECT 1173.5 465.816 1176.5 468.816 ;
        RECT 1243.5 465.816 1246.5 468.816 ;
        RECT 1307.5 465.816 1310.5 468.816 ;
        RECT 1373.5 465.816 1376.5 468.816 ;
        RECT 1443.5 465.816 1446.5 468.816 ;
        RECT 1507.5 465.816 1510.5 468.816 ;
        RECT 1573.5 465.816 1576.5 468.816 ;
    END
  END VSS
  PIN piso_sw_out
    DIRECTION OUTPUT ;
    USE POWER ;
  END piso_sw_out
  PIN sipo_sw_out
    DIRECTION OUTPUT ;
    USE POWER ;
  END sipo_sw_out
  PIN VDDM
    DIRECTION OUTPUT ;
    USE POWER ;
  END VDDM
  OBS
    LAYER M2 ;
      RECT 611.792 467.816 612.92 468.116 ;
      RECT 809.24 467.816 809.912 468.116 ;
      RECT 812.28 465.116 897.768 468.116 ;
      RECT 0.7 0.7 1638.212 468.06 ;
      RECT 899.224 465.116 922.544 468.116 ;
      RECT 924 465.116 1004.928 468.116 ;
      RECT 1006.384 465.116 1197.208 468.116 ;
      RECT 1198.664 465.116 1301.48 468.116 ;
      RECT 1302.936 465.116 1437.52 468.116 ;
      RECT 1438.976 465.116 1486.92 468.116 ;
      RECT 1488.376 465.116 1638.212 468.116 ;
      RECT 0.7 465.116 10.848 468.116 ;
      RECT 12.304 465.116 25.744 468.116 ;
      RECT 27.2 465.116 76.816 468.116 ;
      RECT 78.272 465.116 218.632 468.116 ;
      RECT 220.088 465.116 320.624 468.116 ;
      RECT 322.08 465.116 349.808 468.116 ;
      RECT 351.264 465.116 507.888 468.116 ;
      RECT 509.344 465.116 533.424 468.116 ;
      RECT 534.88 465.116 544.216 468.116 ;
      RECT 545.672 465.116 610.336 468.116 ;
      RECT 614.376 465.116 649.856 468.116 ;
      RECT 651.312 465.116 695.152 468.116 ;
      RECT 696.608 465.116 721.904 468.116 ;
      RECT 723.36 465.116 775.408 468.116 ;
      RECT 776.864 465.116 784.984 468.116 ;
      RECT 786.44 465.116 802.16 468.116 ;
      RECT 803.616 465.116 806.872 468.116 ;
      POLYGON 1335.678 468.695 1335.678 468.585 1335.676 468.585 1335.676 468.116 1437.52 468.116 1437.52 468.06 1438.976 468.06 1438.976 468.116 1486.92 468.116 1486.92 468.06 1488.376 468.06 1488.376 468.116 1638.212 468.116 1638.212 0.7 1613.838 0.7 1613.838 0.577 1613.778 0.577 1613.778 0.7 1612.164 0.7 1612.164 0.403 1612.166 0.403 1612.166 0.273 1612.106 0.273 1612.106 0.403 1612.108 0.403 1612.108 0.7 1204.196 0.7 1204.196 0.403 1204.198 0.403 1204.198 0.273 1204.138 0.273 1204.138 0.403 1204.14 0.403 1204.14 0.7 1173.038 0.7 1173.038 0.577 1172.978 0.577 1172.978 0.7 806.564 0.7 806.564 0.251 806.566 0.251 806.566 0.121 806.506 0.121 806.506 0.251 806.508 0.251 806.508 0.7 694.996 0.7 694.996 0.555 694.998 0.555 694.998 0.425 694.938 0.425 694.938 0.555 694.94 0.555 694.94 0.7 612.31 0.7 612.31 0.577 612.25 0.577 612.25 0.7 49.452 0.7 49.452 0.555 49.454 0.555 49.454 0.425 49.394 0.425 49.394 0.555 49.396 0.555 49.396 0.7 6.742 0.7 6.742 0.577 6.682 0.577 6.682 0.7 5.068 0.7 5.068 0.403 5.07 0.403 5.07 0.273 5.01 0.273 5.01 0.403 5.012 0.403 5.012 0.7 4.004 0.7 4.004 0.251 4.006 0.251 4.006 0.121 3.946 0.121 3.946 0.251 3.948 0.251 3.948 0.7 0.7 0.7 0.7 468.116 10.848 468.116 10.848 468.06 12.304 468.06 12.304 468.116 25.744 468.116 25.744 468.06 27.2 468.06 27.2 468.116 76.816 468.116 76.816 468.06 78.272 468.06 78.272 468.116 218.632 468.116 218.632 468.06 220.088 468.06 220.088 468.116 320.624 468.116 320.624 468.06 322.08 468.06 322.08 468.116 349.808 468.116 349.808 468.06 351.264 468.06 351.264 468.116 507.888 468.116 507.888 468.06 509.344 468.06 509.344 468.116 533.424 468.116 533.424 468.06 534.88 468.06 534.88 468.116 544.216 468.116 544.216 468.06 545.672 468.06 545.672 468.116 610.336 468.116 610.336 468.06 611.792 468.06 611.792 468.116 612.92 468.116 612.92 468.06 614.376 468.06 614.376 468.116 649.856 468.116 649.856 468.06 651.312 468.06 651.312 468.116 695.152 468.116 695.152 468.06 696.608 468.06 696.608 468.116 721.904 468.116 721.904 468.06 723.36 468.06 723.36 468.116 775.408 468.116 775.408 468.06 776.864 468.06 776.864 468.116 784.984 468.116 784.984 468.06 786.44 468.06 786.44 468.116 802.16 468.116 802.16 468.06 803.616 468.06 803.616 468.116 806.872 468.116 806.872 468.06 809.24 468.06 809.24 468.116 809.912 468.116 809.912 468.06 811.068 468.06 811.068 468.565 811.066 468.565 811.066 468.695 811.126 468.695 811.126 468.565 811.124 468.565 811.124 468.06 812.28 468.06 812.28 468.116 897.768 468.116 897.768 468.06 899.224 468.06 899.224 468.116 922.544 468.116 922.544 468.06 924 468.06 924 468.116 1004.928 468.116 1004.928 468.06 1006.384 468.06 1006.384 468.116 1197.208 468.116 1197.208 468.06 1198.664 468.06 1198.664 468.116 1301.48 468.116 1301.48 468.06 1302.936 468.06 1302.936 468.116 1335.62 468.116 1335.62 468.585 1335.618 468.585 1335.618 468.695 ;
      POLYGON 0.206 342.383 0.206 342.253 0.204 342.253 0.204 181.587 0.206 181.587 0.206 181.457 0.146 181.457 0.146 181.587 0.148 181.587 0.148 342.253 0.146 342.253 0.146 342.383 ;
      POLYGON 0.51 337.671 0.51 337.561 0.508 337.561 0.508 180.503 0.51 180.503 0.51 180.393 0.45 180.393 0.45 180.503 0.452 180.503 0.452 337.561 0.45 337.561 0.45 337.671 ;
      POLYGON 0.662 272.007 0.662 271.897 0.66 271.897 0.66 267.143 0.662 267.143 0.662 267.033 0.602 267.033 0.602 267.143 0.604 267.143 0.604 271.897 0.602 271.897 0.602 272.007 ;
      POLYGON 0.662 163.479 0.662 163.349 0.66 163.349 0.66 1.923 0.662 1.923 0.662 1.793 0.602 1.793 0.602 1.923 0.604 1.923 0.604 163.349 0.602 163.349 0.602 163.479 ;
      POLYGON 0.51 157.399 0.51 157.289 0.508 157.289 0.508 3.139 0.51 3.139 0.51 3.009 0.45 3.009 0.45 3.139 0.452 3.139 0.452 157.289 0.45 157.289 0.45 157.399 ;
      POLYGON 0.206 148.735 0.206 148.605 0.204 148.605 0.204 0.251 0.206 0.251 0.206 0.121 0.146 0.121 0.146 0.251 0.148 0.251 0.148 148.605 0.146 148.605 0.146 148.735 ;
      RECT 0.45 2.396 0.51 2.663 ;
    LAYER M8 ;
      RECT 1242.2 465.116 1242.8 468.116 ;
      RECT 1247.2 465.116 1247.8 468.116 ;
      RECT 1306.2 465.116 1306.8 468.116 ;
      RECT 1311.2 465.116 1311.8 468.116 ;
      RECT 1372.2 465.116 1372.8 468.116 ;
      RECT 1377.2 465.116 1377.8 468.116 ;
      RECT 1442.2 465.116 1442.8 468.116 ;
      RECT 1447.2 465.116 1447.8 468.116 ;
      RECT 1506.2 465.116 1506.8 468.116 ;
      RECT 1511.2 465.116 1511.8 468.116 ;
      RECT 1572.2 465.116 1572.8 468.116 ;
      RECT 1577.2 465.116 1577.8 468.116 ;
      RECT 842.2 465.116 842.8 468.116 ;
      RECT 847.2 465.116 847.8 468.116 ;
      RECT 906.2 465.116 906.8 468.116 ;
      RECT 911.2 465.116 911.8 468.116 ;
      RECT 972.2 465.116 972.8 468.116 ;
      RECT 977.2 465.116 977.8 468.116 ;
      RECT 1042.2 465.116 1042.8 468.116 ;
      RECT 1047.2 465.116 1047.8 468.116 ;
      RECT 1106.2 465.116 1106.8 468.116 ;
      RECT 1111.2 465.116 1111.8 468.116 ;
      RECT 1172.2 465.116 1172.8 468.116 ;
      RECT 1177.2 465.116 1177.8 468.116 ;
      RECT 442.2 465.116 442.8 468.116 ;
      RECT 447.2 465.116 447.8 468.116 ;
      RECT 506.2 465.116 506.8 468.116 ;
      RECT 511.2 465.116 511.8 468.116 ;
      RECT 572.2 465.116 572.8 468.116 ;
      RECT 577.2 465.116 577.8 468.116 ;
      RECT 642.2 465.116 642.8 468.116 ;
      RECT 647.2 465.116 647.8 468.116 ;
      RECT 706.2 465.116 706.8 468.116 ;
      RECT 711.2 465.116 711.8 468.116 ;
      RECT 772.2 465.116 772.8 468.116 ;
      RECT 777.2 465.116 777.8 468.116 ;
      RECT 42.2 465.116 42.8 468.116 ;
      RECT 47.2 465.116 47.8 468.116 ;
      RECT 106.2 465.116 106.8 468.116 ;
      RECT 111.2 465.116 111.8 468.116 ;
      RECT 172.2 465.116 172.8 468.116 ;
      RECT 177.2 465.116 177.8 468.116 ;
      RECT 242.2 465.116 242.8 468.116 ;
      RECT 247.2 465.116 247.8 468.116 ;
      RECT 306.2 465.116 306.8 468.116 ;
      RECT 311.2 465.116 311.8 468.116 ;
      RECT 372.2 465.116 372.8 468.116 ;
      RECT 377.2 465.116 377.8 468.116 ;
      RECT 1242.2 0.7 1242.8 3.7 ;
      RECT 1247.2 0.7 1247.8 3.7 ;
      RECT 1306.2 0.7 1306.8 3.7 ;
      RECT 1311.2 0.7 1311.8 3.7 ;
      RECT 1372.2 0.7 1372.8 3.7 ;
      RECT 1377.2 0.7 1377.8 3.7 ;
      RECT 1442.2 0.7 1442.8 3.7 ;
      RECT 1447.2 0.7 1447.8 3.7 ;
      RECT 1506.2 0.7 1506.8 3.7 ;
      RECT 1511.2 0.7 1511.8 3.7 ;
      RECT 1572.2 0.7 1572.8 3.7 ;
      RECT 1577.2 0.7 1577.8 3.7 ;
      RECT 842.2 0.7 842.8 3.7 ;
      RECT 847.2 0.7 847.8 3.7 ;
      RECT 906.2 0.7 906.8 3.7 ;
      RECT 911.2 0.7 911.8 3.7 ;
      RECT 972.2 0.7 972.8 3.7 ;
      RECT 977.2 0.7 977.8 3.7 ;
      RECT 1042.2 0.7 1042.8 3.7 ;
      RECT 1047.2 0.7 1047.8 3.7 ;
      RECT 1106.2 0.7 1106.8 3.7 ;
      RECT 1111.2 0.7 1111.8 3.7 ;
      RECT 1172.2 0.7 1172.8 3.7 ;
      RECT 1177.2 0.7 1177.8 3.7 ;
      RECT 442.2 0.7 442.8 3.7 ;
      RECT 447.2 0.7 447.8 3.7 ;
      RECT 506.2 0.7 506.8 3.7 ;
      RECT 511.2 0.7 511.8 3.7 ;
      RECT 572.2 0.7 572.8 3.7 ;
      RECT 577.2 0.7 577.8 3.7 ;
      RECT 642.2 0.7 642.8 3.7 ;
      RECT 647.2 0.7 647.8 3.7 ;
      RECT 706.2 0.7 706.8 3.7 ;
      RECT 711.2 0.7 711.8 3.7 ;
      RECT 772.2 0.7 772.8 3.7 ;
      RECT 777.2 0.7 777.8 3.7 ;
      RECT 42.2 0.7 42.8 3.7 ;
      RECT 47.2 0.7 47.8 3.7 ;
      RECT 106.2 0.7 106.8 3.7 ;
      RECT 111.2 0.7 111.8 3.7 ;
      RECT 172.2 0.7 172.8 3.7 ;
      RECT 177.2 0.7 177.8 3.7 ;
      RECT 242.2 0.7 242.8 3.7 ;
      RECT 247.2 0.7 247.8 3.7 ;
      RECT 306.2 0.7 306.8 3.7 ;
      RECT 311.2 0.7 311.8 3.7 ;
      RECT 372.2 0.7 372.8 3.7 ;
      RECT 377.2 0.7 377.8 3.7 ;
      RECT 782.2 465.116 837.8 468.116 ;
      RECT 0.7 465.116 37.8 468.116 ;
      RECT 52.2 465.116 101.8 468.116 ;
      RECT 116.2 465.116 167.8 468.116 ;
      RECT 182.2 465.116 237.8 468.116 ;
      RECT 252.2 465.116 301.8 468.116 ;
      RECT 316.2 465.116 367.8 468.116 ;
      RECT 382.2 465.116 437.8 468.116 ;
      RECT 452.2 465.116 501.8 468.116 ;
      RECT 516.2 465.116 567.8 468.116 ;
      RECT 582.2 465.116 637.8 468.116 ;
      RECT 652.2 465.116 701.8 468.116 ;
      RECT 716.2 465.116 767.8 468.116 ;
      RECT 852.2 465.116 901.8 468.116 ;
      RECT 916.2 465.116 967.8 468.116 ;
      RECT 982.2 465.116 1037.8 468.116 ;
      RECT 1052.2 465.116 1101.8 468.116 ;
      RECT 1116.2 465.116 1167.8 468.116 ;
      RECT 1182.2 465.116 1237.8 468.116 ;
      RECT 1252.2 465.116 1301.8 468.116 ;
      RECT 1316.2 465.116 1367.8 468.116 ;
      RECT 1382.2 465.116 1437.8 468.116 ;
      RECT 1452.2 465.116 1501.8 468.116 ;
      RECT 1516.2 465.116 1567.8 468.116 ;
      RECT 1582.2 465.116 1638.212 468.116 ;
      RECT 0.7 3.7 1638.212 465.116 ;
      RECT 782.2 0.7 837.8 3.7 ;
      RECT 852.2 0.7 901.8 3.7 ;
      RECT 916.2 0.7 967.8 3.7 ;
      RECT 982.2 0.7 1037.8 3.7 ;
      RECT 1052.2 0.7 1101.8 3.7 ;
      RECT 1116.2 0.7 1167.8 3.7 ;
      RECT 1182.2 0.7 1237.8 3.7 ;
      RECT 1252.2 0.7 1301.8 3.7 ;
      RECT 1316.2 0.7 1367.8 3.7 ;
      RECT 1382.2 0.7 1437.8 3.7 ;
      RECT 1452.2 0.7 1501.8 3.7 ;
      RECT 1516.2 0.7 1567.8 3.7 ;
      RECT 1582.2 0.7 1638.212 3.7 ;
      RECT 0.7 0.7 37.8 3.7 ;
      RECT 52.2 0.7 101.8 3.7 ;
      RECT 116.2 0.7 167.8 3.7 ;
      RECT 182.2 0.7 237.8 3.7 ;
      RECT 252.2 0.7 301.8 3.7 ;
      RECT 316.2 0.7 367.8 3.7 ;
      RECT 382.2 0.7 437.8 3.7 ;
      RECT 452.2 0.7 501.8 3.7 ;
      RECT 516.2 0.7 567.8 3.7 ;
      RECT 582.2 0.7 637.8 3.7 ;
      RECT 652.2 0.7 701.8 3.7 ;
      RECT 716.2 0.7 767.8 3.7 ;
    LAYER NWELL ;
      RECT 0.23 0.23 1638.682 468.586 ;
    LAYER PO ;
      RECT 0.122 0.122 1638.79 468.694 ;
    LAYER M1 ;
      POLYGON 811.607 468.67 811.607 468.61 811.477 468.61 811.477 468.615 811.171 468.615 811.171 468.61 811.041 468.61 811.041 468.67 811.171 468.67 811.171 468.665 811.477 468.665 811.477 468.67 ;
      RECT 0.75 0.75 1638.162 468.066 ;
      POLYGON 1638.162 468.066 1638.162 0.75 0.75 0.75 0.75 1.823 0.707 1.823 0.707 1.818 0.577 1.818 0.577 1.878 0.707 1.878 0.707 1.873 0.75 1.873 0.75 2.583 0.555 2.583 0.555 2.578 0.425 2.578 0.425 2.638 0.555 2.638 0.555 2.633 0.75 2.633 0.75 3.039 0.555 3.039 0.555 3.034 0.425 3.034 0.425 3.094 0.555 3.094 0.555 3.089 0.75 3.089 0.75 148.655 0.251 148.655 0.251 148.65 0.121 148.65 0.121 148.71 0.251 148.71 0.251 148.705 0.75 148.705 0.75 163.399 0.707 163.399 0.707 163.394 0.577 163.394 0.577 163.454 0.707 163.454 0.707 163.449 0.75 163.449 0.75 181.487 0.251 181.487 0.251 181.482 0.121 181.482 0.121 181.542 0.251 181.542 0.251 181.537 0.75 181.537 0.75 268.426 0.729 268.426 0.729 268.486 0.75 268.486 0.75 342.303 0.251 342.303 0.251 342.298 0.121 342.298 0.121 342.358 0.251 342.358 0.251 342.353 0.75 342.353 0.75 468.066 ;
      POLYGON 1613.863 0.662 1613.863 0.602 1613.733 0.602 1613.733 0.607 1173.083 0.607 1173.083 0.602 1172.953 0.602 1172.953 0.662 1173.083 0.662 1173.083 0.657 1613.733 0.657 1613.733 0.662 ;
      POLYGON 612.335 0.662 612.335 0.602 612.205 0.602 612.205 0.607 6.787 0.607 6.787 0.602 6.657 0.602 6.657 0.662 6.787 0.662 6.787 0.657 612.205 0.657 612.205 0.662 ;
      POLYGON 695.023 0.51 695.023 0.45 694.893 0.45 694.893 0.455 49.499 0.455 49.499 0.45 49.369 0.45 49.369 0.51 49.499 0.51 49.499 0.505 694.893 0.505 694.893 0.51 ;
      POLYGON 1612.191 0.358 1612.191 0.298 1612.061 0.298 1612.061 0.303 1204.243 0.303 1204.243 0.298 1204.113 0.298 1204.113 0.358 1204.243 0.358 1204.243 0.353 1612.061 0.353 1612.061 0.358 ;
      POLYGON 5.095 0.358 5.095 0.298 4.965 0.298 4.965 0.303 4.305 0.303 4.305 0.201 806.461 0.201 806.461 0.206 806.591 0.206 806.591 0.146 806.461 0.146 806.461 0.151 4.255 0.151 4.255 0.353 4.965 0.353 4.965 0.358 ;
      POLYGON 4.031 0.206 4.031 0.146 3.901 0.146 3.901 0.151 0.251 0.151 0.251 0.146 0.121 0.146 0.121 0.206 0.251 0.206 0.251 0.201 3.901 0.201 3.901 0.206 ;
    LAYER VIA1 ;
      RECT 811.527 468.615 811.577 468.665 ;
      RECT 811.071 468.615 811.121 468.665 ;
      RECT 0.151 342.303 0.201 342.353 ;
      RECT 0.151 181.487 0.201 181.537 ;
      RECT 0.607 163.399 0.657 163.449 ;
      RECT 0.151 148.655 0.201 148.705 ;
      RECT 0.455 3.039 0.505 3.089 ;
      RECT 0.455 2.583 0.505 2.633 ;
      RECT 0.607 1.823 0.657 1.873 ;
      RECT 1613.783 0.607 1613.833 0.657 ;
      RECT 1172.983 0.607 1173.033 0.657 ;
      RECT 612.255 0.607 612.305 0.657 ;
      RECT 6.687 0.607 6.737 0.657 ;
      RECT 694.943 0.455 694.993 0.505 ;
      RECT 49.399 0.455 49.449 0.505 ;
      RECT 1612.111 0.303 1612.161 0.353 ;
      RECT 1204.143 0.303 1204.193 0.353 ;
      RECT 5.015 0.303 5.065 0.353 ;
      RECT 806.511 0.151 806.561 0.201 ;
      RECT 3.951 0.151 4.001 0.201 ;
      RECT 0.151 0.151 0.201 0.201 ;
    LAYER VIA2 ;
      RECT 1438.223 468.615 1438.273 468.665 ;
      RECT 1335.623 468.615 1335.673 468.665 ;
      RECT 1197.911 468.615 1197.961 468.665 ;
      RECT 810.919 468.615 810.969 468.665 ;
      RECT 219.335 468.615 219.385 468.665 ;
      RECT 0.455 337.591 0.505 337.641 ;
      RECT 0.607 271.927 0.657 271.977 ;
      RECT 0.607 267.063 0.657 267.113 ;
      RECT 0.455 180.423 0.505 180.473 ;
      RECT 0.455 157.319 0.505 157.369 ;
      RECT 0.455 2.583 0.505 2.633 ;
    LAYER M3 ;
      POLYGON 1438.303 468.67 1438.303 468.61 1438.193 468.61 1438.193 468.612 1335.703 468.612 1335.703 468.61 1335.593 468.61 1335.593 468.67 1335.703 468.67 1335.703 468.668 1438.193 468.668 1438.193 468.67 ;
      POLYGON 1197.991 468.67 1197.991 468.61 1197.881 468.61 1197.881 468.612 1028.359 468.612 1028.359 468.61 1028.249 468.61 1028.249 468.67 1028.359 468.67 1028.359 468.668 1197.881 468.668 1197.881 468.67 ;
      RECT 810.732 468.61 810.999 468.67 ;
      POLYGON 427.351 468.67 427.351 468.61 427.241 468.61 427.241 468.612 219.415 468.612 219.415 468.61 219.305 468.61 219.305 468.67 219.415 468.67 219.415 468.668 427.241 468.668 427.241 468.67 ;
      RECT 0.7 0.7 1638.212 468.116 ;
      POLYGON 1638.212 468.116 1638.212 0.7 406.044 0.7 406.044 0.508 418.604 0.508 418.604 0.7 418.66 0.7 418.66 0.452 405.988 0.452 405.988 0.7 0.7 0.7 0.7 12.916 0.231 12.916 0.231 12.914 0.121 12.914 0.121 12.974 0.231 12.974 0.231 12.972 0.7 12.972 0.7 54.564 0.535 54.564 0.535 54.562 0.425 54.562 0.425 54.622 0.535 54.622 0.535 54.62 0.7 54.62 0.7 54.868 0.535 54.868 0.535 54.866 0.425 54.866 0.425 54.926 0.535 54.926 0.535 54.924 0.7 54.924 0.7 157.316 0.535 157.316 0.535 157.314 0.425 157.314 0.425 157.374 0.535 157.374 0.535 157.372 0.7 157.372 0.7 159.748 0.535 159.748 0.535 159.746 0.425 159.746 0.425 159.806 0.535 159.806 0.535 159.804 0.7 159.804 0.7 175.252 0.231 175.252 0.231 175.25 0.121 175.25 0.121 175.31 0.231 175.31 0.231 175.308 0.7 175.308 0.7 180.42 0.535 180.42 0.535 180.418 0.425 180.418 0.425 180.478 0.535 180.478 0.535 180.476 0.7 180.476 0.7 190.148 0.535 190.148 0.535 190.146 0.425 190.146 0.425 190.206 0.535 190.206 0.535 190.204 0.7 190.204 0.7 265.54 0.231 265.54 0.231 265.538 0.121 265.538 0.121 265.598 0.231 265.598 0.231 265.596 0.7 265.596 0.7 266.148 0.231 266.148 0.231 266.146 0.121 266.146 0.121 266.206 0.231 266.206 0.231 266.204 0.7 266.204 0.7 267.97 0.572 267.97 0.572 268.03 0.7 268.03 0.7 271.924 0.687 271.924 0.687 271.922 0.577 271.922 0.577 271.982 0.687 271.982 0.687 271.98 0.7 271.98 0.7 293.508 0.231 293.508 0.231 293.506 0.121 293.506 0.121 293.566 0.231 293.566 0.231 293.564 0.7 293.564 0.7 294.724 0.231 294.724 0.231 294.722 0.121 294.722 0.121 294.782 0.231 294.782 0.231 294.78 0.7 294.78 0.7 336.068 0.231 336.068 0.231 336.066 0.121 336.066 0.121 336.126 0.231 336.126 0.231 336.124 0.7 336.124 0.7 337.588 0.535 337.588 0.535 337.586 0.425 337.586 0.425 337.646 0.535 337.646 0.535 337.644 0.7 337.644 0.7 468.116 ;
      RECT 0.42 267.058 0.687 267.118 ;
      RECT 0.268 2.578 0.535 2.638 ;
      POLYGON 1613.863 0.51 1613.863 0.45 1613.753 0.45 1613.753 0.452 1407.143 0.452 1407.143 0.45 1407.033 0.45 1407.033 0.51 1407.143 0.51 1407.143 0.508 1613.753 0.508 1613.753 0.51 ;
      POLYGON 405.463 0.206 405.463 0.146 405.353 0.146 405.353 0.148 196.615 0.148 196.615 0.146 196.505 0.146 196.505 0.206 196.615 0.206 196.615 0.204 405.353 0.204 405.353 0.206 ;
      POLYGON 172.295 0.206 172.295 0.146 172.185 0.146 172.185 0.148 2.967 0.148 2.967 0.146 2.857 0.146 2.857 0.206 2.967 0.206 2.967 0.204 172.185 0.204 172.185 0.206 ;
    LAYER VIA3 ;
      RECT 1028.279 468.615 1028.329 468.665 ;
      RECT 810.919 468.615 810.969 468.665 ;
      RECT 427.271 468.615 427.321 468.665 ;
      RECT 0.151 336.071 0.201 336.121 ;
      RECT 0.151 294.727 0.201 294.777 ;
      RECT 0.151 293.511 0.201 293.561 ;
      RECT 0.607 267.063 0.657 267.113 ;
      RECT 0.151 266.151 0.201 266.201 ;
      RECT 0.151 265.543 0.201 265.593 ;
      RECT 0.455 190.151 0.505 190.201 ;
      RECT 0.151 175.255 0.201 175.305 ;
      RECT 0.455 159.751 0.505 159.801 ;
      RECT 0.455 54.871 0.505 54.921 ;
      RECT 0.455 54.567 0.505 54.617 ;
      RECT 0.151 12.919 0.201 12.969 ;
      RECT 0.455 2.583 0.505 2.633 ;
      RECT 1613.783 0.455 1613.833 0.505 ;
      RECT 1407.063 0.455 1407.113 0.505 ;
      RECT 405.383 0.151 405.433 0.201 ;
      RECT 196.535 0.151 196.585 0.201 ;
      RECT 172.215 0.151 172.265 0.201 ;
      RECT 2.887 0.151 2.937 0.201 ;
    LAYER M4 ;
      RECT 0.7 0.7 1638.212 468.116 ;
      POLYGON 1028.334 468.695 1028.334 468.585 1028.332 468.585 1028.332 468.116 1638.212 468.116 1638.212 0.7 1618.396 0.7 1618.396 0.231 1618.398 0.231 1618.398 0.121 1618.338 0.121 1618.338 0.231 1618.34 0.231 1618.34 0.7 1613.836 0.7 1613.836 0.535 1613.838 0.535 1613.838 0.425 1613.778 0.425 1613.778 0.535 1613.78 0.535 1613.78 0.7 1407.116 0.7 1407.116 0.535 1407.118 0.535 1407.118 0.425 1407.058 0.425 1407.058 0.535 1407.06 0.535 1407.06 0.7 405.436 0.7 405.436 0.231 405.438 0.231 405.438 0.121 405.378 0.121 405.378 0.231 405.38 0.231 405.38 0.7 213.918 0.7 213.918 0.572 213.858 0.572 213.858 0.7 213.612 0.7 213.612 0.231 213.614 0.231 213.614 0.121 213.554 0.121 213.554 0.231 213.556 0.231 213.556 0.7 206.62 0.7 206.62 0.231 206.622 0.231 206.622 0.121 206.562 0.121 206.562 0.231 206.564 0.231 206.564 0.7 196.588 0.7 196.588 0.231 196.59 0.231 196.59 0.121 196.53 0.121 196.53 0.231 196.532 0.231 196.532 0.7 172.268 0.7 172.268 0.231 172.27 0.231 172.27 0.121 172.21 0.121 172.21 0.231 172.212 0.231 172.212 0.7 54.316 0.7 54.316 0.231 54.318 0.231 54.318 0.121 54.258 0.121 54.258 0.231 54.26 0.231 54.26 0.7 50.972 0.7 50.972 0.231 50.974 0.231 50.974 0.121 50.914 0.121 50.914 0.231 50.916 0.231 50.916 0.7 34.252 0.7 34.252 0.231 34.254 0.231 34.254 0.121 34.194 0.121 34.194 0.231 34.196 0.231 34.196 0.7 6.588 0.7 6.588 0.231 6.59 0.231 6.59 0.121 6.53 0.121 6.53 0.231 6.532 0.231 6.532 0.7 2.94 0.7 2.94 0.231 2.942 0.231 2.942 0.121 2.882 0.121 2.882 0.231 2.884 0.231 2.884 0.7 0.7 0.7 0.7 468.116 427.268 468.116 427.268 468.585 427.266 468.585 427.266 468.695 427.326 468.695 427.326 468.585 427.324 468.585 427.324 468.116 810.916 468.116 810.916 468.585 810.914 468.585 810.914 468.695 810.974 468.695 810.974 468.585 810.972 468.585 810.972 468.116 1028.276 468.116 1028.276 468.585 1028.274 468.585 1028.274 468.695 ;
      POLYGON 0.206 336.151 0.206 336.041 0.204 336.041 0.204 294.807 0.206 294.807 0.206 294.697 0.146 294.697 0.146 294.807 0.148 294.807 0.148 336.041 0.146 336.041 0.146 336.151 ;
      POLYGON 0.51 334.023 0.51 333.913 0.508 333.913 0.508 190.231 0.51 190.231 0.51 190.121 0.45 190.121 0.45 190.231 0.452 190.231 0.452 333.913 0.45 333.913 0.45 334.023 ;
      POLYGON 0.206 293.591 0.206 293.481 0.204 293.481 0.204 266.231 0.206 266.231 0.206 266.121 0.146 266.121 0.146 266.231 0.148 266.231 0.148 293.481 0.146 293.481 0.146 293.591 ;
      RECT 0.602 266.876 0.662 267.143 ;
      POLYGON 0.206 265.623 0.206 265.513 0.204 265.513 0.204 175.335 0.206 175.335 0.206 175.225 0.146 175.225 0.146 175.335 0.148 175.335 0.148 265.513 0.146 265.513 0.146 265.623 ;
      POLYGON 0.51 159.831 0.51 159.721 0.508 159.721 0.508 54.951 0.51 54.951 0.51 54.841 0.45 54.841 0.45 54.951 0.452 54.951 0.452 159.721 0.45 159.721 0.45 159.831 ;
      POLYGON 0.206 127.911 0.206 127.801 0.204 127.801 0.204 12.999 0.206 12.999 0.206 12.889 0.146 12.889 0.146 12.999 0.148 12.999 0.148 127.801 0.146 127.801 0.146 127.911 ;
      POLYGON 0.51 54.647 0.51 54.537 0.508 54.537 0.508 2.663 0.51 2.663 0.51 2.553 0.45 2.553 0.45 2.663 0.452 2.663 0.452 54.537 0.45 54.537 0.45 54.647 ;
    LAYER VIA4 ;
      RECT 0.455 333.943 0.505 333.993 ;
      RECT 0.607 267.063 0.657 267.113 ;
      RECT 0.151 127.831 0.201 127.881 ;
      RECT 1618.343 0.151 1618.393 0.201 ;
      RECT 213.559 0.151 213.609 0.201 ;
      RECT 206.567 0.151 206.617 0.201 ;
      RECT 54.263 0.151 54.313 0.201 ;
      RECT 50.919 0.151 50.969 0.201 ;
      RECT 34.199 0.151 34.249 0.201 ;
      RECT 6.535 0.151 6.585 0.201 ;
    LAYER M5 ;
      RECT 0.7 0.7 1638.212 468.116 ;
      POLYGON 1638.212 468.116 1638.212 0.7 32.732 0.7 32.732 0.148 6.615 0.148 6.615 0.146 6.505 0.146 6.505 0.206 6.615 0.206 6.615 0.204 32.676 0.204 32.676 0.7 0.7 0.7 0.7 3.188 0.231 3.188 0.231 3.186 0.121 3.186 0.121 3.246 0.231 3.246 0.231 3.244 0.7 3.244 0.7 108.978 0.572 108.978 0.572 109.038 0.7 109.038 0.7 112.02 0.231 112.02 0.231 112.018 0.121 112.018 0.121 112.078 0.231 112.078 0.231 112.076 0.7 112.076 0.7 113.844 0.231 113.844 0.231 113.842 0.121 113.842 0.121 113.902 0.231 113.902 0.231 113.9 0.7 113.9 0.7 127.828 0.231 127.828 0.231 127.826 0.121 127.826 0.121 127.886 0.231 127.886 0.231 127.884 0.7 127.884 0.7 158.228 0.231 158.228 0.231 158.226 0.121 158.226 0.121 158.286 0.231 158.286 0.231 158.284 0.7 158.284 0.7 190.45 0.572 190.45 0.572 190.51 0.7 190.51 0.7 191.668 0.231 191.668 0.231 191.666 0.121 191.666 0.121 191.726 0.231 191.726 0.231 191.724 0.7 191.724 0.7 268.276 0.231 268.276 0.231 268.274 0.121 268.274 0.121 268.334 0.231 268.334 0.231 268.332 0.7 268.332 0.7 333.94 0.535 333.94 0.535 333.938 0.425 333.938 0.425 333.998 0.535 333.998 0.535 333.996 0.7 333.996 0.7 358.868 0.231 358.868 0.231 358.866 0.121 358.866 0.121 358.926 0.231 358.926 0.231 358.924 0.7 358.924 0.7 468.116 ;
      POLYGON 0.687 267.118 0.687 267.058 0.577 267.058 0.577 267.06 0.231 267.06 0.231 267.058 0.121 267.058 0.121 267.118 0.231 267.118 0.231 267.116 0.577 267.116 0.577 267.118 ;
      POLYGON 1618.423 0.206 1618.423 0.146 1618.313 0.146 1618.313 0.148 1408.359 0.148 1408.359 0.146 1408.249 0.146 1408.249 0.206 1408.359 0.206 1408.359 0.204 1618.313 0.204 1618.313 0.206 ;
      POLYGON 555.335 0.206 555.335 0.146 555.225 0.146 555.225 0.148 213.639 0.148 213.639 0.146 213.529 0.146 213.529 0.206 213.639 0.206 213.639 0.204 555.225 0.204 555.225 0.206 ;
      POLYGON 206.647 0.206 206.647 0.146 206.537 0.146 206.537 0.148 54.343 0.148 54.343 0.146 54.233 0.146 54.233 0.206 54.343 0.206 54.343 0.204 206.537 0.204 206.537 0.206 ;
      POLYGON 50.999 0.206 50.999 0.146 50.889 0.146 50.889 0.148 34.279 0.148 34.279 0.146 34.169 0.146 34.169 0.206 34.279 0.206 34.279 0.204 50.889 0.204 50.889 0.206 ;
    LAYER VIA5 ;
      RECT 0.151 358.871 0.201 358.921 ;
      RECT 0.151 268.279 0.201 268.329 ;
      RECT 0.151 267.063 0.201 267.113 ;
      RECT 0.151 191.671 0.201 191.721 ;
      RECT 0.151 158.231 0.201 158.281 ;
      RECT 0.151 113.847 0.201 113.897 ;
      RECT 0.151 112.023 0.201 112.073 ;
      RECT 0.151 3.191 0.201 3.241 ;
      RECT 1408.279 0.151 1408.329 0.201 ;
      RECT 555.255 0.151 555.305 0.201 ;
    LAYER M6 ;
      RECT 0.7 0.7 1638.212 468.116 ;
      POLYGON 1638.212 468.116 1638.212 0.7 1408.332 0.7 1408.332 0.231 1408.334 0.231 1408.334 0.121 1408.274 0.121 1408.274 0.231 1408.276 0.231 1408.276 0.7 555.308 0.7 555.308 0.231 555.31 0.231 555.31 0.121 555.25 0.121 555.25 0.231 555.252 0.231 555.252 0.7 0.7 0.7 0.7 468.116 ;
      POLYGON 0.206 358.951 0.206 358.841 0.204 358.841 0.204 268.359 0.206 268.359 0.206 268.249 0.146 268.249 0.146 268.359 0.148 268.359 0.148 358.841 0.146 358.841 0.146 358.951 ;
      POLYGON 0.206 267.143 0.206 267.033 0.204 267.033 0.204 191.751 0.206 191.751 0.206 191.641 0.146 191.641 0.146 191.751 0.148 191.751 0.148 267.033 0.146 267.033 0.146 267.143 ;
      POLYGON 0.206 158.311 0.206 158.201 0.204 158.201 0.204 113.927 0.206 113.927 0.206 113.817 0.146 113.817 0.146 113.927 0.148 113.927 0.148 158.201 0.146 158.201 0.146 158.311 ;
      POLYGON 0.206 112.103 0.206 111.993 0.204 111.993 0.204 3.271 0.206 3.271 0.206 3.161 0.146 3.161 0.146 3.271 0.148 3.271 0.148 111.993 0.146 111.993 0.146 112.103 ;
    LAYER M7 ;
      RECT 0.7 0.7 1638.212 468.116 ;
    LAYER VIA7 ;
      RECT 1571.415 466.791 1571.465 466.841 ;
      RECT 1571.295 466.791 1571.345 466.841 ;
      RECT 1571.175 466.791 1571.225 466.841 ;
      RECT 1571.055 466.791 1571.105 466.841 ;
      RECT 1570.935 466.791 1570.985 466.841 ;
      RECT 1570.815 466.791 1570.865 466.841 ;
      RECT 1570.695 466.791 1570.745 466.841 ;
      RECT 1570.575 466.791 1570.625 466.841 ;
      RECT 1570.455 466.791 1570.505 466.841 ;
      RECT 1570.335 466.791 1570.385 466.841 ;
      RECT 1570.215 466.791 1570.265 466.841 ;
      RECT 1570.095 466.791 1570.145 466.841 ;
      RECT 1569.975 466.791 1570.025 466.841 ;
      RECT 1569.855 466.791 1569.905 466.841 ;
      RECT 1569.735 466.791 1569.785 466.841 ;
      RECT 1569.615 466.791 1569.665 466.841 ;
      RECT 1569.495 466.791 1569.545 466.841 ;
      RECT 1569.375 466.791 1569.425 466.841 ;
      RECT 1569.255 466.791 1569.305 466.841 ;
      RECT 1569.135 466.791 1569.185 466.841 ;
      RECT 1569.015 466.791 1569.065 466.841 ;
      RECT 1568.895 466.791 1568.945 466.841 ;
      RECT 1568.775 466.791 1568.825 466.841 ;
      RECT 1568.655 466.791 1568.705 466.841 ;
      RECT 1568.535 466.791 1568.585 466.841 ;
      RECT 1505.415 466.791 1505.465 466.841 ;
      RECT 1505.295 466.791 1505.345 466.841 ;
      RECT 1505.175 466.791 1505.225 466.841 ;
      RECT 1505.055 466.791 1505.105 466.841 ;
      RECT 1504.935 466.791 1504.985 466.841 ;
      RECT 1504.815 466.791 1504.865 466.841 ;
      RECT 1504.695 466.791 1504.745 466.841 ;
      RECT 1504.575 466.791 1504.625 466.841 ;
      RECT 1504.455 466.791 1504.505 466.841 ;
      RECT 1504.335 466.791 1504.385 466.841 ;
      RECT 1504.215 466.791 1504.265 466.841 ;
      RECT 1504.095 466.791 1504.145 466.841 ;
      RECT 1503.975 466.791 1504.025 466.841 ;
      RECT 1503.855 466.791 1503.905 466.841 ;
      RECT 1503.735 466.791 1503.785 466.841 ;
      RECT 1503.615 466.791 1503.665 466.841 ;
      RECT 1503.495 466.791 1503.545 466.841 ;
      RECT 1503.375 466.791 1503.425 466.841 ;
      RECT 1503.255 466.791 1503.305 466.841 ;
      RECT 1503.135 466.791 1503.185 466.841 ;
      RECT 1503.015 466.791 1503.065 466.841 ;
      RECT 1502.895 466.791 1502.945 466.841 ;
      RECT 1502.775 466.791 1502.825 466.841 ;
      RECT 1502.655 466.791 1502.705 466.841 ;
      RECT 1502.535 466.791 1502.585 466.841 ;
      RECT 1441.415 466.791 1441.465 466.841 ;
      RECT 1441.295 466.791 1441.345 466.841 ;
      RECT 1441.175 466.791 1441.225 466.841 ;
      RECT 1441.055 466.791 1441.105 466.841 ;
      RECT 1440.935 466.791 1440.985 466.841 ;
      RECT 1440.815 466.791 1440.865 466.841 ;
      RECT 1440.695 466.791 1440.745 466.841 ;
      RECT 1440.575 466.791 1440.625 466.841 ;
      RECT 1440.455 466.791 1440.505 466.841 ;
      RECT 1440.335 466.791 1440.385 466.841 ;
      RECT 1440.215 466.791 1440.265 466.841 ;
      RECT 1440.095 466.791 1440.145 466.841 ;
      RECT 1439.975 466.791 1440.025 466.841 ;
      RECT 1439.855 466.791 1439.905 466.841 ;
      RECT 1439.735 466.791 1439.785 466.841 ;
      RECT 1439.615 466.791 1439.665 466.841 ;
      RECT 1439.495 466.791 1439.545 466.841 ;
      RECT 1439.375 466.791 1439.425 466.841 ;
      RECT 1439.255 466.791 1439.305 466.841 ;
      RECT 1439.135 466.791 1439.185 466.841 ;
      RECT 1439.015 466.791 1439.065 466.841 ;
      RECT 1438.895 466.791 1438.945 466.841 ;
      RECT 1438.775 466.791 1438.825 466.841 ;
      RECT 1438.655 466.791 1438.705 466.841 ;
      RECT 1438.535 466.791 1438.585 466.841 ;
      RECT 1371.415 466.791 1371.465 466.841 ;
      RECT 1371.295 466.791 1371.345 466.841 ;
      RECT 1371.175 466.791 1371.225 466.841 ;
      RECT 1371.055 466.791 1371.105 466.841 ;
      RECT 1370.935 466.791 1370.985 466.841 ;
      RECT 1370.815 466.791 1370.865 466.841 ;
      RECT 1370.695 466.791 1370.745 466.841 ;
      RECT 1370.575 466.791 1370.625 466.841 ;
      RECT 1370.455 466.791 1370.505 466.841 ;
      RECT 1370.335 466.791 1370.385 466.841 ;
      RECT 1370.215 466.791 1370.265 466.841 ;
      RECT 1370.095 466.791 1370.145 466.841 ;
      RECT 1369.975 466.791 1370.025 466.841 ;
      RECT 1369.855 466.791 1369.905 466.841 ;
      RECT 1369.735 466.791 1369.785 466.841 ;
      RECT 1369.615 466.791 1369.665 466.841 ;
      RECT 1369.495 466.791 1369.545 466.841 ;
      RECT 1369.375 466.791 1369.425 466.841 ;
      RECT 1369.255 466.791 1369.305 466.841 ;
      RECT 1369.135 466.791 1369.185 466.841 ;
      RECT 1369.015 466.791 1369.065 466.841 ;
      RECT 1368.895 466.791 1368.945 466.841 ;
      RECT 1368.775 466.791 1368.825 466.841 ;
      RECT 1368.655 466.791 1368.705 466.841 ;
      RECT 1368.535 466.791 1368.585 466.841 ;
      RECT 1305.415 466.791 1305.465 466.841 ;
      RECT 1305.295 466.791 1305.345 466.841 ;
      RECT 1305.175 466.791 1305.225 466.841 ;
      RECT 1305.055 466.791 1305.105 466.841 ;
      RECT 1304.935 466.791 1304.985 466.841 ;
      RECT 1304.815 466.791 1304.865 466.841 ;
      RECT 1304.695 466.791 1304.745 466.841 ;
      RECT 1304.575 466.791 1304.625 466.841 ;
      RECT 1304.455 466.791 1304.505 466.841 ;
      RECT 1304.335 466.791 1304.385 466.841 ;
      RECT 1304.215 466.791 1304.265 466.841 ;
      RECT 1304.095 466.791 1304.145 466.841 ;
      RECT 1303.975 466.791 1304.025 466.841 ;
      RECT 1303.855 466.791 1303.905 466.841 ;
      RECT 1303.735 466.791 1303.785 466.841 ;
      RECT 1303.615 466.791 1303.665 466.841 ;
      RECT 1303.495 466.791 1303.545 466.841 ;
      RECT 1303.375 466.791 1303.425 466.841 ;
      RECT 1303.255 466.791 1303.305 466.841 ;
      RECT 1303.135 466.791 1303.185 466.841 ;
      RECT 1303.015 466.791 1303.065 466.841 ;
      RECT 1302.895 466.791 1302.945 466.841 ;
      RECT 1302.775 466.791 1302.825 466.841 ;
      RECT 1302.655 466.791 1302.705 466.841 ;
      RECT 1302.535 466.791 1302.585 466.841 ;
      RECT 1241.415 466.791 1241.465 466.841 ;
      RECT 1241.295 466.791 1241.345 466.841 ;
      RECT 1241.175 466.791 1241.225 466.841 ;
      RECT 1241.055 466.791 1241.105 466.841 ;
      RECT 1240.935 466.791 1240.985 466.841 ;
      RECT 1240.815 466.791 1240.865 466.841 ;
      RECT 1240.695 466.791 1240.745 466.841 ;
      RECT 1240.575 466.791 1240.625 466.841 ;
      RECT 1240.455 466.791 1240.505 466.841 ;
      RECT 1240.335 466.791 1240.385 466.841 ;
      RECT 1240.215 466.791 1240.265 466.841 ;
      RECT 1240.095 466.791 1240.145 466.841 ;
      RECT 1239.975 466.791 1240.025 466.841 ;
      RECT 1239.855 466.791 1239.905 466.841 ;
      RECT 1239.735 466.791 1239.785 466.841 ;
      RECT 1239.615 466.791 1239.665 466.841 ;
      RECT 1239.495 466.791 1239.545 466.841 ;
      RECT 1239.375 466.791 1239.425 466.841 ;
      RECT 1239.255 466.791 1239.305 466.841 ;
      RECT 1239.135 466.791 1239.185 466.841 ;
      RECT 1239.015 466.791 1239.065 466.841 ;
      RECT 1238.895 466.791 1238.945 466.841 ;
      RECT 1238.775 466.791 1238.825 466.841 ;
      RECT 1238.655 466.791 1238.705 466.841 ;
      RECT 1238.535 466.791 1238.585 466.841 ;
      RECT 1171.415 466.791 1171.465 466.841 ;
      RECT 1171.295 466.791 1171.345 466.841 ;
      RECT 1171.175 466.791 1171.225 466.841 ;
      RECT 1171.055 466.791 1171.105 466.841 ;
      RECT 1170.935 466.791 1170.985 466.841 ;
      RECT 1170.815 466.791 1170.865 466.841 ;
      RECT 1170.695 466.791 1170.745 466.841 ;
      RECT 1170.575 466.791 1170.625 466.841 ;
      RECT 1170.455 466.791 1170.505 466.841 ;
      RECT 1170.335 466.791 1170.385 466.841 ;
      RECT 1170.215 466.791 1170.265 466.841 ;
      RECT 1170.095 466.791 1170.145 466.841 ;
      RECT 1169.975 466.791 1170.025 466.841 ;
      RECT 1169.855 466.791 1169.905 466.841 ;
      RECT 1169.735 466.791 1169.785 466.841 ;
      RECT 1169.615 466.791 1169.665 466.841 ;
      RECT 1169.495 466.791 1169.545 466.841 ;
      RECT 1169.375 466.791 1169.425 466.841 ;
      RECT 1169.255 466.791 1169.305 466.841 ;
      RECT 1169.135 466.791 1169.185 466.841 ;
      RECT 1169.015 466.791 1169.065 466.841 ;
      RECT 1168.895 466.791 1168.945 466.841 ;
      RECT 1168.775 466.791 1168.825 466.841 ;
      RECT 1168.655 466.791 1168.705 466.841 ;
      RECT 1168.535 466.791 1168.585 466.841 ;
      RECT 1105.415 466.791 1105.465 466.841 ;
      RECT 1105.295 466.791 1105.345 466.841 ;
      RECT 1105.175 466.791 1105.225 466.841 ;
      RECT 1105.055 466.791 1105.105 466.841 ;
      RECT 1104.935 466.791 1104.985 466.841 ;
      RECT 1104.815 466.791 1104.865 466.841 ;
      RECT 1104.695 466.791 1104.745 466.841 ;
      RECT 1104.575 466.791 1104.625 466.841 ;
      RECT 1104.455 466.791 1104.505 466.841 ;
      RECT 1104.335 466.791 1104.385 466.841 ;
      RECT 1104.215 466.791 1104.265 466.841 ;
      RECT 1104.095 466.791 1104.145 466.841 ;
      RECT 1103.975 466.791 1104.025 466.841 ;
      RECT 1103.855 466.791 1103.905 466.841 ;
      RECT 1103.735 466.791 1103.785 466.841 ;
      RECT 1103.615 466.791 1103.665 466.841 ;
      RECT 1103.495 466.791 1103.545 466.841 ;
      RECT 1103.375 466.791 1103.425 466.841 ;
      RECT 1103.255 466.791 1103.305 466.841 ;
      RECT 1103.135 466.791 1103.185 466.841 ;
      RECT 1103.015 466.791 1103.065 466.841 ;
      RECT 1102.895 466.791 1102.945 466.841 ;
      RECT 1102.775 466.791 1102.825 466.841 ;
      RECT 1102.655 466.791 1102.705 466.841 ;
      RECT 1102.535 466.791 1102.585 466.841 ;
      RECT 1041.415 466.791 1041.465 466.841 ;
      RECT 1041.295 466.791 1041.345 466.841 ;
      RECT 1041.175 466.791 1041.225 466.841 ;
      RECT 1041.055 466.791 1041.105 466.841 ;
      RECT 1040.935 466.791 1040.985 466.841 ;
      RECT 1040.815 466.791 1040.865 466.841 ;
      RECT 1040.695 466.791 1040.745 466.841 ;
      RECT 1040.575 466.791 1040.625 466.841 ;
      RECT 1040.455 466.791 1040.505 466.841 ;
      RECT 1040.335 466.791 1040.385 466.841 ;
      RECT 1040.215 466.791 1040.265 466.841 ;
      RECT 1040.095 466.791 1040.145 466.841 ;
      RECT 1039.975 466.791 1040.025 466.841 ;
      RECT 1039.855 466.791 1039.905 466.841 ;
      RECT 1039.735 466.791 1039.785 466.841 ;
      RECT 1039.615 466.791 1039.665 466.841 ;
      RECT 1039.495 466.791 1039.545 466.841 ;
      RECT 1039.375 466.791 1039.425 466.841 ;
      RECT 1039.255 466.791 1039.305 466.841 ;
      RECT 1039.135 466.791 1039.185 466.841 ;
      RECT 1039.015 466.791 1039.065 466.841 ;
      RECT 1038.895 466.791 1038.945 466.841 ;
      RECT 1038.775 466.791 1038.825 466.841 ;
      RECT 1038.655 466.791 1038.705 466.841 ;
      RECT 1038.535 466.791 1038.585 466.841 ;
      RECT 971.415 466.791 971.465 466.841 ;
      RECT 971.295 466.791 971.345 466.841 ;
      RECT 971.175 466.791 971.225 466.841 ;
      RECT 971.055 466.791 971.105 466.841 ;
      RECT 970.935 466.791 970.985 466.841 ;
      RECT 970.815 466.791 970.865 466.841 ;
      RECT 970.695 466.791 970.745 466.841 ;
      RECT 970.575 466.791 970.625 466.841 ;
      RECT 970.455 466.791 970.505 466.841 ;
      RECT 970.335 466.791 970.385 466.841 ;
      RECT 970.215 466.791 970.265 466.841 ;
      RECT 970.095 466.791 970.145 466.841 ;
      RECT 969.975 466.791 970.025 466.841 ;
      RECT 969.855 466.791 969.905 466.841 ;
      RECT 969.735 466.791 969.785 466.841 ;
      RECT 969.615 466.791 969.665 466.841 ;
      RECT 969.495 466.791 969.545 466.841 ;
      RECT 969.375 466.791 969.425 466.841 ;
      RECT 969.255 466.791 969.305 466.841 ;
      RECT 969.135 466.791 969.185 466.841 ;
      RECT 969.015 466.791 969.065 466.841 ;
      RECT 968.895 466.791 968.945 466.841 ;
      RECT 968.775 466.791 968.825 466.841 ;
      RECT 968.655 466.791 968.705 466.841 ;
      RECT 968.535 466.791 968.585 466.841 ;
      RECT 905.415 466.791 905.465 466.841 ;
      RECT 905.295 466.791 905.345 466.841 ;
      RECT 905.175 466.791 905.225 466.841 ;
      RECT 905.055 466.791 905.105 466.841 ;
      RECT 904.935 466.791 904.985 466.841 ;
      RECT 904.815 466.791 904.865 466.841 ;
      RECT 904.695 466.791 904.745 466.841 ;
      RECT 904.575 466.791 904.625 466.841 ;
      RECT 904.455 466.791 904.505 466.841 ;
      RECT 904.335 466.791 904.385 466.841 ;
      RECT 904.215 466.791 904.265 466.841 ;
      RECT 904.095 466.791 904.145 466.841 ;
      RECT 903.975 466.791 904.025 466.841 ;
      RECT 903.855 466.791 903.905 466.841 ;
      RECT 903.735 466.791 903.785 466.841 ;
      RECT 903.615 466.791 903.665 466.841 ;
      RECT 903.495 466.791 903.545 466.841 ;
      RECT 903.375 466.791 903.425 466.841 ;
      RECT 903.255 466.791 903.305 466.841 ;
      RECT 903.135 466.791 903.185 466.841 ;
      RECT 903.015 466.791 903.065 466.841 ;
      RECT 902.895 466.791 902.945 466.841 ;
      RECT 902.775 466.791 902.825 466.841 ;
      RECT 902.655 466.791 902.705 466.841 ;
      RECT 902.535 466.791 902.585 466.841 ;
      RECT 841.415 466.791 841.465 466.841 ;
      RECT 841.295 466.791 841.345 466.841 ;
      RECT 841.175 466.791 841.225 466.841 ;
      RECT 841.055 466.791 841.105 466.841 ;
      RECT 840.935 466.791 840.985 466.841 ;
      RECT 840.815 466.791 840.865 466.841 ;
      RECT 840.695 466.791 840.745 466.841 ;
      RECT 840.575 466.791 840.625 466.841 ;
      RECT 840.455 466.791 840.505 466.841 ;
      RECT 840.335 466.791 840.385 466.841 ;
      RECT 840.215 466.791 840.265 466.841 ;
      RECT 840.095 466.791 840.145 466.841 ;
      RECT 839.975 466.791 840.025 466.841 ;
      RECT 839.855 466.791 839.905 466.841 ;
      RECT 839.735 466.791 839.785 466.841 ;
      RECT 839.615 466.791 839.665 466.841 ;
      RECT 839.495 466.791 839.545 466.841 ;
      RECT 839.375 466.791 839.425 466.841 ;
      RECT 839.255 466.791 839.305 466.841 ;
      RECT 839.135 466.791 839.185 466.841 ;
      RECT 839.015 466.791 839.065 466.841 ;
      RECT 838.895 466.791 838.945 466.841 ;
      RECT 838.775 466.791 838.825 466.841 ;
      RECT 838.655 466.791 838.705 466.841 ;
      RECT 838.535 466.791 838.585 466.841 ;
      RECT 771.415 466.791 771.465 466.841 ;
      RECT 771.295 466.791 771.345 466.841 ;
      RECT 771.175 466.791 771.225 466.841 ;
      RECT 771.055 466.791 771.105 466.841 ;
      RECT 770.935 466.791 770.985 466.841 ;
      RECT 770.815 466.791 770.865 466.841 ;
      RECT 770.695 466.791 770.745 466.841 ;
      RECT 770.575 466.791 770.625 466.841 ;
      RECT 770.455 466.791 770.505 466.841 ;
      RECT 770.335 466.791 770.385 466.841 ;
      RECT 770.215 466.791 770.265 466.841 ;
      RECT 770.095 466.791 770.145 466.841 ;
      RECT 769.975 466.791 770.025 466.841 ;
      RECT 769.855 466.791 769.905 466.841 ;
      RECT 769.735 466.791 769.785 466.841 ;
      RECT 769.615 466.791 769.665 466.841 ;
      RECT 769.495 466.791 769.545 466.841 ;
      RECT 769.375 466.791 769.425 466.841 ;
      RECT 769.255 466.791 769.305 466.841 ;
      RECT 769.135 466.791 769.185 466.841 ;
      RECT 769.015 466.791 769.065 466.841 ;
      RECT 768.895 466.791 768.945 466.841 ;
      RECT 768.775 466.791 768.825 466.841 ;
      RECT 768.655 466.791 768.705 466.841 ;
      RECT 768.535 466.791 768.585 466.841 ;
      RECT 705.415 466.791 705.465 466.841 ;
      RECT 705.295 466.791 705.345 466.841 ;
      RECT 705.175 466.791 705.225 466.841 ;
      RECT 705.055 466.791 705.105 466.841 ;
      RECT 704.935 466.791 704.985 466.841 ;
      RECT 704.815 466.791 704.865 466.841 ;
      RECT 704.695 466.791 704.745 466.841 ;
      RECT 704.575 466.791 704.625 466.841 ;
      RECT 704.455 466.791 704.505 466.841 ;
      RECT 704.335 466.791 704.385 466.841 ;
      RECT 704.215 466.791 704.265 466.841 ;
      RECT 704.095 466.791 704.145 466.841 ;
      RECT 703.975 466.791 704.025 466.841 ;
      RECT 703.855 466.791 703.905 466.841 ;
      RECT 703.735 466.791 703.785 466.841 ;
      RECT 703.615 466.791 703.665 466.841 ;
      RECT 703.495 466.791 703.545 466.841 ;
      RECT 703.375 466.791 703.425 466.841 ;
      RECT 703.255 466.791 703.305 466.841 ;
      RECT 703.135 466.791 703.185 466.841 ;
      RECT 703.015 466.791 703.065 466.841 ;
      RECT 702.895 466.791 702.945 466.841 ;
      RECT 702.775 466.791 702.825 466.841 ;
      RECT 702.655 466.791 702.705 466.841 ;
      RECT 702.535 466.791 702.585 466.841 ;
      RECT 641.415 466.791 641.465 466.841 ;
      RECT 641.295 466.791 641.345 466.841 ;
      RECT 641.175 466.791 641.225 466.841 ;
      RECT 641.055 466.791 641.105 466.841 ;
      RECT 640.935 466.791 640.985 466.841 ;
      RECT 640.815 466.791 640.865 466.841 ;
      RECT 640.695 466.791 640.745 466.841 ;
      RECT 640.575 466.791 640.625 466.841 ;
      RECT 640.455 466.791 640.505 466.841 ;
      RECT 640.335 466.791 640.385 466.841 ;
      RECT 640.215 466.791 640.265 466.841 ;
      RECT 640.095 466.791 640.145 466.841 ;
      RECT 639.975 466.791 640.025 466.841 ;
      RECT 639.855 466.791 639.905 466.841 ;
      RECT 639.735 466.791 639.785 466.841 ;
      RECT 639.615 466.791 639.665 466.841 ;
      RECT 639.495 466.791 639.545 466.841 ;
      RECT 639.375 466.791 639.425 466.841 ;
      RECT 639.255 466.791 639.305 466.841 ;
      RECT 639.135 466.791 639.185 466.841 ;
      RECT 639.015 466.791 639.065 466.841 ;
      RECT 638.895 466.791 638.945 466.841 ;
      RECT 638.775 466.791 638.825 466.841 ;
      RECT 638.655 466.791 638.705 466.841 ;
      RECT 638.535 466.791 638.585 466.841 ;
      RECT 571.415 466.791 571.465 466.841 ;
      RECT 571.295 466.791 571.345 466.841 ;
      RECT 571.175 466.791 571.225 466.841 ;
      RECT 571.055 466.791 571.105 466.841 ;
      RECT 570.935 466.791 570.985 466.841 ;
      RECT 570.815 466.791 570.865 466.841 ;
      RECT 570.695 466.791 570.745 466.841 ;
      RECT 570.575 466.791 570.625 466.841 ;
      RECT 570.455 466.791 570.505 466.841 ;
      RECT 570.335 466.791 570.385 466.841 ;
      RECT 570.215 466.791 570.265 466.841 ;
      RECT 570.095 466.791 570.145 466.841 ;
      RECT 569.975 466.791 570.025 466.841 ;
      RECT 569.855 466.791 569.905 466.841 ;
      RECT 569.735 466.791 569.785 466.841 ;
      RECT 569.615 466.791 569.665 466.841 ;
      RECT 569.495 466.791 569.545 466.841 ;
      RECT 569.375 466.791 569.425 466.841 ;
      RECT 569.255 466.791 569.305 466.841 ;
      RECT 569.135 466.791 569.185 466.841 ;
      RECT 569.015 466.791 569.065 466.841 ;
      RECT 568.895 466.791 568.945 466.841 ;
      RECT 568.775 466.791 568.825 466.841 ;
      RECT 568.655 466.791 568.705 466.841 ;
      RECT 568.535 466.791 568.585 466.841 ;
      RECT 505.415 466.791 505.465 466.841 ;
      RECT 505.295 466.791 505.345 466.841 ;
      RECT 505.175 466.791 505.225 466.841 ;
      RECT 505.055 466.791 505.105 466.841 ;
      RECT 504.935 466.791 504.985 466.841 ;
      RECT 504.815 466.791 504.865 466.841 ;
      RECT 504.695 466.791 504.745 466.841 ;
      RECT 504.575 466.791 504.625 466.841 ;
      RECT 504.455 466.791 504.505 466.841 ;
      RECT 504.335 466.791 504.385 466.841 ;
      RECT 504.215 466.791 504.265 466.841 ;
      RECT 504.095 466.791 504.145 466.841 ;
      RECT 503.975 466.791 504.025 466.841 ;
      RECT 503.855 466.791 503.905 466.841 ;
      RECT 503.735 466.791 503.785 466.841 ;
      RECT 503.615 466.791 503.665 466.841 ;
      RECT 503.495 466.791 503.545 466.841 ;
      RECT 503.375 466.791 503.425 466.841 ;
      RECT 503.255 466.791 503.305 466.841 ;
      RECT 503.135 466.791 503.185 466.841 ;
      RECT 503.015 466.791 503.065 466.841 ;
      RECT 502.895 466.791 502.945 466.841 ;
      RECT 502.775 466.791 502.825 466.841 ;
      RECT 502.655 466.791 502.705 466.841 ;
      RECT 502.535 466.791 502.585 466.841 ;
      RECT 441.415 466.791 441.465 466.841 ;
      RECT 441.295 466.791 441.345 466.841 ;
      RECT 441.175 466.791 441.225 466.841 ;
      RECT 441.055 466.791 441.105 466.841 ;
      RECT 440.935 466.791 440.985 466.841 ;
      RECT 440.815 466.791 440.865 466.841 ;
      RECT 440.695 466.791 440.745 466.841 ;
      RECT 440.575 466.791 440.625 466.841 ;
      RECT 440.455 466.791 440.505 466.841 ;
      RECT 440.335 466.791 440.385 466.841 ;
      RECT 440.215 466.791 440.265 466.841 ;
      RECT 440.095 466.791 440.145 466.841 ;
      RECT 439.975 466.791 440.025 466.841 ;
      RECT 439.855 466.791 439.905 466.841 ;
      RECT 439.735 466.791 439.785 466.841 ;
      RECT 439.615 466.791 439.665 466.841 ;
      RECT 439.495 466.791 439.545 466.841 ;
      RECT 439.375 466.791 439.425 466.841 ;
      RECT 439.255 466.791 439.305 466.841 ;
      RECT 439.135 466.791 439.185 466.841 ;
      RECT 439.015 466.791 439.065 466.841 ;
      RECT 438.895 466.791 438.945 466.841 ;
      RECT 438.775 466.791 438.825 466.841 ;
      RECT 438.655 466.791 438.705 466.841 ;
      RECT 438.535 466.791 438.585 466.841 ;
      RECT 371.415 466.791 371.465 466.841 ;
      RECT 371.295 466.791 371.345 466.841 ;
      RECT 371.175 466.791 371.225 466.841 ;
      RECT 371.055 466.791 371.105 466.841 ;
      RECT 370.935 466.791 370.985 466.841 ;
      RECT 370.815 466.791 370.865 466.841 ;
      RECT 370.695 466.791 370.745 466.841 ;
      RECT 370.575 466.791 370.625 466.841 ;
      RECT 370.455 466.791 370.505 466.841 ;
      RECT 370.335 466.791 370.385 466.841 ;
      RECT 370.215 466.791 370.265 466.841 ;
      RECT 370.095 466.791 370.145 466.841 ;
      RECT 369.975 466.791 370.025 466.841 ;
      RECT 369.855 466.791 369.905 466.841 ;
      RECT 369.735 466.791 369.785 466.841 ;
      RECT 369.615 466.791 369.665 466.841 ;
      RECT 369.495 466.791 369.545 466.841 ;
      RECT 369.375 466.791 369.425 466.841 ;
      RECT 369.255 466.791 369.305 466.841 ;
      RECT 369.135 466.791 369.185 466.841 ;
      RECT 369.015 466.791 369.065 466.841 ;
      RECT 368.895 466.791 368.945 466.841 ;
      RECT 368.775 466.791 368.825 466.841 ;
      RECT 368.655 466.791 368.705 466.841 ;
      RECT 368.535 466.791 368.585 466.841 ;
      RECT 305.415 466.791 305.465 466.841 ;
      RECT 305.295 466.791 305.345 466.841 ;
      RECT 305.175 466.791 305.225 466.841 ;
      RECT 305.055 466.791 305.105 466.841 ;
      RECT 304.935 466.791 304.985 466.841 ;
      RECT 304.815 466.791 304.865 466.841 ;
      RECT 304.695 466.791 304.745 466.841 ;
      RECT 304.575 466.791 304.625 466.841 ;
      RECT 304.455 466.791 304.505 466.841 ;
      RECT 304.335 466.791 304.385 466.841 ;
      RECT 304.215 466.791 304.265 466.841 ;
      RECT 304.095 466.791 304.145 466.841 ;
      RECT 303.975 466.791 304.025 466.841 ;
      RECT 303.855 466.791 303.905 466.841 ;
      RECT 303.735 466.791 303.785 466.841 ;
      RECT 303.615 466.791 303.665 466.841 ;
      RECT 303.495 466.791 303.545 466.841 ;
      RECT 303.375 466.791 303.425 466.841 ;
      RECT 303.255 466.791 303.305 466.841 ;
      RECT 303.135 466.791 303.185 466.841 ;
      RECT 303.015 466.791 303.065 466.841 ;
      RECT 302.895 466.791 302.945 466.841 ;
      RECT 302.775 466.791 302.825 466.841 ;
      RECT 302.655 466.791 302.705 466.841 ;
      RECT 302.535 466.791 302.585 466.841 ;
      RECT 241.415 466.791 241.465 466.841 ;
      RECT 241.295 466.791 241.345 466.841 ;
      RECT 241.175 466.791 241.225 466.841 ;
      RECT 241.055 466.791 241.105 466.841 ;
      RECT 240.935 466.791 240.985 466.841 ;
      RECT 240.815 466.791 240.865 466.841 ;
      RECT 240.695 466.791 240.745 466.841 ;
      RECT 240.575 466.791 240.625 466.841 ;
      RECT 240.455 466.791 240.505 466.841 ;
      RECT 240.335 466.791 240.385 466.841 ;
      RECT 240.215 466.791 240.265 466.841 ;
      RECT 240.095 466.791 240.145 466.841 ;
      RECT 239.975 466.791 240.025 466.841 ;
      RECT 239.855 466.791 239.905 466.841 ;
      RECT 239.735 466.791 239.785 466.841 ;
      RECT 239.615 466.791 239.665 466.841 ;
      RECT 239.495 466.791 239.545 466.841 ;
      RECT 239.375 466.791 239.425 466.841 ;
      RECT 239.255 466.791 239.305 466.841 ;
      RECT 239.135 466.791 239.185 466.841 ;
      RECT 239.015 466.791 239.065 466.841 ;
      RECT 238.895 466.791 238.945 466.841 ;
      RECT 238.775 466.791 238.825 466.841 ;
      RECT 238.655 466.791 238.705 466.841 ;
      RECT 238.535 466.791 238.585 466.841 ;
      RECT 171.415 466.791 171.465 466.841 ;
      RECT 171.295 466.791 171.345 466.841 ;
      RECT 171.175 466.791 171.225 466.841 ;
      RECT 171.055 466.791 171.105 466.841 ;
      RECT 170.935 466.791 170.985 466.841 ;
      RECT 170.815 466.791 170.865 466.841 ;
      RECT 170.695 466.791 170.745 466.841 ;
      RECT 170.575 466.791 170.625 466.841 ;
      RECT 170.455 466.791 170.505 466.841 ;
      RECT 170.335 466.791 170.385 466.841 ;
      RECT 170.215 466.791 170.265 466.841 ;
      RECT 170.095 466.791 170.145 466.841 ;
      RECT 169.975 466.791 170.025 466.841 ;
      RECT 169.855 466.791 169.905 466.841 ;
      RECT 169.735 466.791 169.785 466.841 ;
      RECT 169.615 466.791 169.665 466.841 ;
      RECT 169.495 466.791 169.545 466.841 ;
      RECT 169.375 466.791 169.425 466.841 ;
      RECT 169.255 466.791 169.305 466.841 ;
      RECT 169.135 466.791 169.185 466.841 ;
      RECT 169.015 466.791 169.065 466.841 ;
      RECT 168.895 466.791 168.945 466.841 ;
      RECT 168.775 466.791 168.825 466.841 ;
      RECT 168.655 466.791 168.705 466.841 ;
      RECT 168.535 466.791 168.585 466.841 ;
      RECT 105.415 466.791 105.465 466.841 ;
      RECT 105.295 466.791 105.345 466.841 ;
      RECT 105.175 466.791 105.225 466.841 ;
      RECT 105.055 466.791 105.105 466.841 ;
      RECT 104.935 466.791 104.985 466.841 ;
      RECT 104.815 466.791 104.865 466.841 ;
      RECT 104.695 466.791 104.745 466.841 ;
      RECT 104.575 466.791 104.625 466.841 ;
      RECT 104.455 466.791 104.505 466.841 ;
      RECT 104.335 466.791 104.385 466.841 ;
      RECT 104.215 466.791 104.265 466.841 ;
      RECT 104.095 466.791 104.145 466.841 ;
      RECT 103.975 466.791 104.025 466.841 ;
      RECT 103.855 466.791 103.905 466.841 ;
      RECT 103.735 466.791 103.785 466.841 ;
      RECT 103.615 466.791 103.665 466.841 ;
      RECT 103.495 466.791 103.545 466.841 ;
      RECT 103.375 466.791 103.425 466.841 ;
      RECT 103.255 466.791 103.305 466.841 ;
      RECT 103.135 466.791 103.185 466.841 ;
      RECT 103.015 466.791 103.065 466.841 ;
      RECT 102.895 466.791 102.945 466.841 ;
      RECT 102.775 466.791 102.825 466.841 ;
      RECT 102.655 466.791 102.705 466.841 ;
      RECT 102.535 466.791 102.585 466.841 ;
      RECT 41.415 466.791 41.465 466.841 ;
      RECT 41.295 466.791 41.345 466.841 ;
      RECT 41.175 466.791 41.225 466.841 ;
      RECT 41.055 466.791 41.105 466.841 ;
      RECT 40.935 466.791 40.985 466.841 ;
      RECT 40.815 466.791 40.865 466.841 ;
      RECT 40.695 466.791 40.745 466.841 ;
      RECT 40.575 466.791 40.625 466.841 ;
      RECT 40.455 466.791 40.505 466.841 ;
      RECT 40.335 466.791 40.385 466.841 ;
      RECT 40.215 466.791 40.265 466.841 ;
      RECT 40.095 466.791 40.145 466.841 ;
      RECT 39.975 466.791 40.025 466.841 ;
      RECT 39.855 466.791 39.905 466.841 ;
      RECT 39.735 466.791 39.785 466.841 ;
      RECT 39.615 466.791 39.665 466.841 ;
      RECT 39.495 466.791 39.545 466.841 ;
      RECT 39.375 466.791 39.425 466.841 ;
      RECT 39.255 466.791 39.305 466.841 ;
      RECT 39.135 466.791 39.185 466.841 ;
      RECT 39.015 466.791 39.065 466.841 ;
      RECT 38.895 466.791 38.945 466.841 ;
      RECT 38.775 466.791 38.825 466.841 ;
      RECT 38.655 466.791 38.705 466.841 ;
      RECT 38.535 466.791 38.585 466.841 ;
      RECT 1576.415 465.119 1576.465 465.169 ;
      RECT 1576.295 465.119 1576.345 465.169 ;
      RECT 1576.175 465.119 1576.225 465.169 ;
      RECT 1576.055 465.119 1576.105 465.169 ;
      RECT 1575.935 465.119 1575.985 465.169 ;
      RECT 1575.815 465.119 1575.865 465.169 ;
      RECT 1575.695 465.119 1575.745 465.169 ;
      RECT 1575.575 465.119 1575.625 465.169 ;
      RECT 1575.455 465.119 1575.505 465.169 ;
      RECT 1575.335 465.119 1575.385 465.169 ;
      RECT 1575.215 465.119 1575.265 465.169 ;
      RECT 1575.095 465.119 1575.145 465.169 ;
      RECT 1574.975 465.119 1575.025 465.169 ;
      RECT 1574.855 465.119 1574.905 465.169 ;
      RECT 1574.735 465.119 1574.785 465.169 ;
      RECT 1574.615 465.119 1574.665 465.169 ;
      RECT 1574.495 465.119 1574.545 465.169 ;
      RECT 1574.375 465.119 1574.425 465.169 ;
      RECT 1574.255 465.119 1574.305 465.169 ;
      RECT 1574.135 465.119 1574.185 465.169 ;
      RECT 1574.015 465.119 1574.065 465.169 ;
      RECT 1573.895 465.119 1573.945 465.169 ;
      RECT 1573.775 465.119 1573.825 465.169 ;
      RECT 1573.655 465.119 1573.705 465.169 ;
      RECT 1573.535 465.119 1573.585 465.169 ;
      RECT 1510.415 465.119 1510.465 465.169 ;
      RECT 1510.295 465.119 1510.345 465.169 ;
      RECT 1510.175 465.119 1510.225 465.169 ;
      RECT 1510.055 465.119 1510.105 465.169 ;
      RECT 1509.935 465.119 1509.985 465.169 ;
      RECT 1509.815 465.119 1509.865 465.169 ;
      RECT 1509.695 465.119 1509.745 465.169 ;
      RECT 1509.575 465.119 1509.625 465.169 ;
      RECT 1509.455 465.119 1509.505 465.169 ;
      RECT 1509.335 465.119 1509.385 465.169 ;
      RECT 1509.215 465.119 1509.265 465.169 ;
      RECT 1509.095 465.119 1509.145 465.169 ;
      RECT 1508.975 465.119 1509.025 465.169 ;
      RECT 1508.855 465.119 1508.905 465.169 ;
      RECT 1508.735 465.119 1508.785 465.169 ;
      RECT 1508.615 465.119 1508.665 465.169 ;
      RECT 1508.495 465.119 1508.545 465.169 ;
      RECT 1508.375 465.119 1508.425 465.169 ;
      RECT 1508.255 465.119 1508.305 465.169 ;
      RECT 1508.135 465.119 1508.185 465.169 ;
      RECT 1508.015 465.119 1508.065 465.169 ;
      RECT 1507.895 465.119 1507.945 465.169 ;
      RECT 1507.775 465.119 1507.825 465.169 ;
      RECT 1507.655 465.119 1507.705 465.169 ;
      RECT 1507.535 465.119 1507.585 465.169 ;
      RECT 1446.415 465.119 1446.465 465.169 ;
      RECT 1446.295 465.119 1446.345 465.169 ;
      RECT 1446.175 465.119 1446.225 465.169 ;
      RECT 1446.055 465.119 1446.105 465.169 ;
      RECT 1445.935 465.119 1445.985 465.169 ;
      RECT 1445.815 465.119 1445.865 465.169 ;
      RECT 1445.695 465.119 1445.745 465.169 ;
      RECT 1445.575 465.119 1445.625 465.169 ;
      RECT 1445.455 465.119 1445.505 465.169 ;
      RECT 1445.335 465.119 1445.385 465.169 ;
      RECT 1445.215 465.119 1445.265 465.169 ;
      RECT 1445.095 465.119 1445.145 465.169 ;
      RECT 1444.975 465.119 1445.025 465.169 ;
      RECT 1444.855 465.119 1444.905 465.169 ;
      RECT 1444.735 465.119 1444.785 465.169 ;
      RECT 1444.615 465.119 1444.665 465.169 ;
      RECT 1444.495 465.119 1444.545 465.169 ;
      RECT 1444.375 465.119 1444.425 465.169 ;
      RECT 1444.255 465.119 1444.305 465.169 ;
      RECT 1444.135 465.119 1444.185 465.169 ;
      RECT 1444.015 465.119 1444.065 465.169 ;
      RECT 1443.895 465.119 1443.945 465.169 ;
      RECT 1443.775 465.119 1443.825 465.169 ;
      RECT 1443.655 465.119 1443.705 465.169 ;
      RECT 1443.535 465.119 1443.585 465.169 ;
      RECT 1376.415 465.119 1376.465 465.169 ;
      RECT 1376.295 465.119 1376.345 465.169 ;
      RECT 1376.175 465.119 1376.225 465.169 ;
      RECT 1376.055 465.119 1376.105 465.169 ;
      RECT 1375.935 465.119 1375.985 465.169 ;
      RECT 1375.815 465.119 1375.865 465.169 ;
      RECT 1375.695 465.119 1375.745 465.169 ;
      RECT 1375.575 465.119 1375.625 465.169 ;
      RECT 1375.455 465.119 1375.505 465.169 ;
      RECT 1375.335 465.119 1375.385 465.169 ;
      RECT 1375.215 465.119 1375.265 465.169 ;
      RECT 1375.095 465.119 1375.145 465.169 ;
      RECT 1374.975 465.119 1375.025 465.169 ;
      RECT 1374.855 465.119 1374.905 465.169 ;
      RECT 1374.735 465.119 1374.785 465.169 ;
      RECT 1374.615 465.119 1374.665 465.169 ;
      RECT 1374.495 465.119 1374.545 465.169 ;
      RECT 1374.375 465.119 1374.425 465.169 ;
      RECT 1374.255 465.119 1374.305 465.169 ;
      RECT 1374.135 465.119 1374.185 465.169 ;
      RECT 1374.015 465.119 1374.065 465.169 ;
      RECT 1373.895 465.119 1373.945 465.169 ;
      RECT 1373.775 465.119 1373.825 465.169 ;
      RECT 1373.655 465.119 1373.705 465.169 ;
      RECT 1373.535 465.119 1373.585 465.169 ;
      RECT 1310.415 465.119 1310.465 465.169 ;
      RECT 1310.295 465.119 1310.345 465.169 ;
      RECT 1310.175 465.119 1310.225 465.169 ;
      RECT 1310.055 465.119 1310.105 465.169 ;
      RECT 1309.935 465.119 1309.985 465.169 ;
      RECT 1309.815 465.119 1309.865 465.169 ;
      RECT 1309.695 465.119 1309.745 465.169 ;
      RECT 1309.575 465.119 1309.625 465.169 ;
      RECT 1309.455 465.119 1309.505 465.169 ;
      RECT 1309.335 465.119 1309.385 465.169 ;
      RECT 1309.215 465.119 1309.265 465.169 ;
      RECT 1309.095 465.119 1309.145 465.169 ;
      RECT 1308.975 465.119 1309.025 465.169 ;
      RECT 1308.855 465.119 1308.905 465.169 ;
      RECT 1308.735 465.119 1308.785 465.169 ;
      RECT 1308.615 465.119 1308.665 465.169 ;
      RECT 1308.495 465.119 1308.545 465.169 ;
      RECT 1308.375 465.119 1308.425 465.169 ;
      RECT 1308.255 465.119 1308.305 465.169 ;
      RECT 1308.135 465.119 1308.185 465.169 ;
      RECT 1308.015 465.119 1308.065 465.169 ;
      RECT 1307.895 465.119 1307.945 465.169 ;
      RECT 1307.775 465.119 1307.825 465.169 ;
      RECT 1307.655 465.119 1307.705 465.169 ;
      RECT 1307.535 465.119 1307.585 465.169 ;
      RECT 1246.415 465.119 1246.465 465.169 ;
      RECT 1246.295 465.119 1246.345 465.169 ;
      RECT 1246.175 465.119 1246.225 465.169 ;
      RECT 1246.055 465.119 1246.105 465.169 ;
      RECT 1245.935 465.119 1245.985 465.169 ;
      RECT 1245.815 465.119 1245.865 465.169 ;
      RECT 1245.695 465.119 1245.745 465.169 ;
      RECT 1245.575 465.119 1245.625 465.169 ;
      RECT 1245.455 465.119 1245.505 465.169 ;
      RECT 1245.335 465.119 1245.385 465.169 ;
      RECT 1245.215 465.119 1245.265 465.169 ;
      RECT 1245.095 465.119 1245.145 465.169 ;
      RECT 1244.975 465.119 1245.025 465.169 ;
      RECT 1244.855 465.119 1244.905 465.169 ;
      RECT 1244.735 465.119 1244.785 465.169 ;
      RECT 1244.615 465.119 1244.665 465.169 ;
      RECT 1244.495 465.119 1244.545 465.169 ;
      RECT 1244.375 465.119 1244.425 465.169 ;
      RECT 1244.255 465.119 1244.305 465.169 ;
      RECT 1244.135 465.119 1244.185 465.169 ;
      RECT 1244.015 465.119 1244.065 465.169 ;
      RECT 1243.895 465.119 1243.945 465.169 ;
      RECT 1243.775 465.119 1243.825 465.169 ;
      RECT 1243.655 465.119 1243.705 465.169 ;
      RECT 1243.535 465.119 1243.585 465.169 ;
      RECT 1176.415 465.119 1176.465 465.169 ;
      RECT 1176.295 465.119 1176.345 465.169 ;
      RECT 1176.175 465.119 1176.225 465.169 ;
      RECT 1176.055 465.119 1176.105 465.169 ;
      RECT 1175.935 465.119 1175.985 465.169 ;
      RECT 1175.815 465.119 1175.865 465.169 ;
      RECT 1175.695 465.119 1175.745 465.169 ;
      RECT 1175.575 465.119 1175.625 465.169 ;
      RECT 1175.455 465.119 1175.505 465.169 ;
      RECT 1175.335 465.119 1175.385 465.169 ;
      RECT 1175.215 465.119 1175.265 465.169 ;
      RECT 1175.095 465.119 1175.145 465.169 ;
      RECT 1174.975 465.119 1175.025 465.169 ;
      RECT 1174.855 465.119 1174.905 465.169 ;
      RECT 1174.735 465.119 1174.785 465.169 ;
      RECT 1174.615 465.119 1174.665 465.169 ;
      RECT 1174.495 465.119 1174.545 465.169 ;
      RECT 1174.375 465.119 1174.425 465.169 ;
      RECT 1174.255 465.119 1174.305 465.169 ;
      RECT 1174.135 465.119 1174.185 465.169 ;
      RECT 1174.015 465.119 1174.065 465.169 ;
      RECT 1173.895 465.119 1173.945 465.169 ;
      RECT 1173.775 465.119 1173.825 465.169 ;
      RECT 1173.655 465.119 1173.705 465.169 ;
      RECT 1173.535 465.119 1173.585 465.169 ;
      RECT 1110.415 465.119 1110.465 465.169 ;
      RECT 1110.295 465.119 1110.345 465.169 ;
      RECT 1110.175 465.119 1110.225 465.169 ;
      RECT 1110.055 465.119 1110.105 465.169 ;
      RECT 1109.935 465.119 1109.985 465.169 ;
      RECT 1109.815 465.119 1109.865 465.169 ;
      RECT 1109.695 465.119 1109.745 465.169 ;
      RECT 1109.575 465.119 1109.625 465.169 ;
      RECT 1109.455 465.119 1109.505 465.169 ;
      RECT 1109.335 465.119 1109.385 465.169 ;
      RECT 1109.215 465.119 1109.265 465.169 ;
      RECT 1109.095 465.119 1109.145 465.169 ;
      RECT 1108.975 465.119 1109.025 465.169 ;
      RECT 1108.855 465.119 1108.905 465.169 ;
      RECT 1108.735 465.119 1108.785 465.169 ;
      RECT 1108.615 465.119 1108.665 465.169 ;
      RECT 1108.495 465.119 1108.545 465.169 ;
      RECT 1108.375 465.119 1108.425 465.169 ;
      RECT 1108.255 465.119 1108.305 465.169 ;
      RECT 1108.135 465.119 1108.185 465.169 ;
      RECT 1108.015 465.119 1108.065 465.169 ;
      RECT 1107.895 465.119 1107.945 465.169 ;
      RECT 1107.775 465.119 1107.825 465.169 ;
      RECT 1107.655 465.119 1107.705 465.169 ;
      RECT 1107.535 465.119 1107.585 465.169 ;
      RECT 1046.415 465.119 1046.465 465.169 ;
      RECT 1046.295 465.119 1046.345 465.169 ;
      RECT 1046.175 465.119 1046.225 465.169 ;
      RECT 1046.055 465.119 1046.105 465.169 ;
      RECT 1045.935 465.119 1045.985 465.169 ;
      RECT 1045.815 465.119 1045.865 465.169 ;
      RECT 1045.695 465.119 1045.745 465.169 ;
      RECT 1045.575 465.119 1045.625 465.169 ;
      RECT 1045.455 465.119 1045.505 465.169 ;
      RECT 1045.335 465.119 1045.385 465.169 ;
      RECT 1045.215 465.119 1045.265 465.169 ;
      RECT 1045.095 465.119 1045.145 465.169 ;
      RECT 1044.975 465.119 1045.025 465.169 ;
      RECT 1044.855 465.119 1044.905 465.169 ;
      RECT 1044.735 465.119 1044.785 465.169 ;
      RECT 1044.615 465.119 1044.665 465.169 ;
      RECT 1044.495 465.119 1044.545 465.169 ;
      RECT 1044.375 465.119 1044.425 465.169 ;
      RECT 1044.255 465.119 1044.305 465.169 ;
      RECT 1044.135 465.119 1044.185 465.169 ;
      RECT 1044.015 465.119 1044.065 465.169 ;
      RECT 1043.895 465.119 1043.945 465.169 ;
      RECT 1043.775 465.119 1043.825 465.169 ;
      RECT 1043.655 465.119 1043.705 465.169 ;
      RECT 1043.535 465.119 1043.585 465.169 ;
      RECT 976.415 465.119 976.465 465.169 ;
      RECT 976.295 465.119 976.345 465.169 ;
      RECT 976.175 465.119 976.225 465.169 ;
      RECT 976.055 465.119 976.105 465.169 ;
      RECT 975.935 465.119 975.985 465.169 ;
      RECT 975.815 465.119 975.865 465.169 ;
      RECT 975.695 465.119 975.745 465.169 ;
      RECT 975.575 465.119 975.625 465.169 ;
      RECT 975.455 465.119 975.505 465.169 ;
      RECT 975.335 465.119 975.385 465.169 ;
      RECT 975.215 465.119 975.265 465.169 ;
      RECT 975.095 465.119 975.145 465.169 ;
      RECT 974.975 465.119 975.025 465.169 ;
      RECT 974.855 465.119 974.905 465.169 ;
      RECT 974.735 465.119 974.785 465.169 ;
      RECT 974.615 465.119 974.665 465.169 ;
      RECT 974.495 465.119 974.545 465.169 ;
      RECT 974.375 465.119 974.425 465.169 ;
      RECT 974.255 465.119 974.305 465.169 ;
      RECT 974.135 465.119 974.185 465.169 ;
      RECT 974.015 465.119 974.065 465.169 ;
      RECT 973.895 465.119 973.945 465.169 ;
      RECT 973.775 465.119 973.825 465.169 ;
      RECT 973.655 465.119 973.705 465.169 ;
      RECT 973.535 465.119 973.585 465.169 ;
      RECT 910.415 465.119 910.465 465.169 ;
      RECT 910.295 465.119 910.345 465.169 ;
      RECT 910.175 465.119 910.225 465.169 ;
      RECT 910.055 465.119 910.105 465.169 ;
      RECT 909.935 465.119 909.985 465.169 ;
      RECT 909.815 465.119 909.865 465.169 ;
      RECT 909.695 465.119 909.745 465.169 ;
      RECT 909.575 465.119 909.625 465.169 ;
      RECT 909.455 465.119 909.505 465.169 ;
      RECT 909.335 465.119 909.385 465.169 ;
      RECT 909.215 465.119 909.265 465.169 ;
      RECT 909.095 465.119 909.145 465.169 ;
      RECT 908.975 465.119 909.025 465.169 ;
      RECT 908.855 465.119 908.905 465.169 ;
      RECT 908.735 465.119 908.785 465.169 ;
      RECT 908.615 465.119 908.665 465.169 ;
      RECT 908.495 465.119 908.545 465.169 ;
      RECT 908.375 465.119 908.425 465.169 ;
      RECT 908.255 465.119 908.305 465.169 ;
      RECT 908.135 465.119 908.185 465.169 ;
      RECT 908.015 465.119 908.065 465.169 ;
      RECT 907.895 465.119 907.945 465.169 ;
      RECT 907.775 465.119 907.825 465.169 ;
      RECT 907.655 465.119 907.705 465.169 ;
      RECT 907.535 465.119 907.585 465.169 ;
      RECT 846.415 465.119 846.465 465.169 ;
      RECT 846.295 465.119 846.345 465.169 ;
      RECT 846.175 465.119 846.225 465.169 ;
      RECT 846.055 465.119 846.105 465.169 ;
      RECT 845.935 465.119 845.985 465.169 ;
      RECT 845.815 465.119 845.865 465.169 ;
      RECT 845.695 465.119 845.745 465.169 ;
      RECT 845.575 465.119 845.625 465.169 ;
      RECT 845.455 465.119 845.505 465.169 ;
      RECT 845.335 465.119 845.385 465.169 ;
      RECT 845.215 465.119 845.265 465.169 ;
      RECT 845.095 465.119 845.145 465.169 ;
      RECT 844.975 465.119 845.025 465.169 ;
      RECT 844.855 465.119 844.905 465.169 ;
      RECT 844.735 465.119 844.785 465.169 ;
      RECT 844.615 465.119 844.665 465.169 ;
      RECT 844.495 465.119 844.545 465.169 ;
      RECT 844.375 465.119 844.425 465.169 ;
      RECT 844.255 465.119 844.305 465.169 ;
      RECT 844.135 465.119 844.185 465.169 ;
      RECT 844.015 465.119 844.065 465.169 ;
      RECT 843.895 465.119 843.945 465.169 ;
      RECT 843.775 465.119 843.825 465.169 ;
      RECT 843.655 465.119 843.705 465.169 ;
      RECT 843.535 465.119 843.585 465.169 ;
      RECT 776.415 465.119 776.465 465.169 ;
      RECT 776.295 465.119 776.345 465.169 ;
      RECT 776.175 465.119 776.225 465.169 ;
      RECT 776.055 465.119 776.105 465.169 ;
      RECT 775.935 465.119 775.985 465.169 ;
      RECT 775.815 465.119 775.865 465.169 ;
      RECT 775.695 465.119 775.745 465.169 ;
      RECT 775.575 465.119 775.625 465.169 ;
      RECT 775.455 465.119 775.505 465.169 ;
      RECT 775.335 465.119 775.385 465.169 ;
      RECT 775.215 465.119 775.265 465.169 ;
      RECT 775.095 465.119 775.145 465.169 ;
      RECT 774.975 465.119 775.025 465.169 ;
      RECT 774.855 465.119 774.905 465.169 ;
      RECT 774.735 465.119 774.785 465.169 ;
      RECT 774.615 465.119 774.665 465.169 ;
      RECT 774.495 465.119 774.545 465.169 ;
      RECT 774.375 465.119 774.425 465.169 ;
      RECT 774.255 465.119 774.305 465.169 ;
      RECT 774.135 465.119 774.185 465.169 ;
      RECT 774.015 465.119 774.065 465.169 ;
      RECT 773.895 465.119 773.945 465.169 ;
      RECT 773.775 465.119 773.825 465.169 ;
      RECT 773.655 465.119 773.705 465.169 ;
      RECT 773.535 465.119 773.585 465.169 ;
      RECT 710.415 465.119 710.465 465.169 ;
      RECT 710.295 465.119 710.345 465.169 ;
      RECT 710.175 465.119 710.225 465.169 ;
      RECT 710.055 465.119 710.105 465.169 ;
      RECT 709.935 465.119 709.985 465.169 ;
      RECT 709.815 465.119 709.865 465.169 ;
      RECT 709.695 465.119 709.745 465.169 ;
      RECT 709.575 465.119 709.625 465.169 ;
      RECT 709.455 465.119 709.505 465.169 ;
      RECT 709.335 465.119 709.385 465.169 ;
      RECT 709.215 465.119 709.265 465.169 ;
      RECT 709.095 465.119 709.145 465.169 ;
      RECT 708.975 465.119 709.025 465.169 ;
      RECT 708.855 465.119 708.905 465.169 ;
      RECT 708.735 465.119 708.785 465.169 ;
      RECT 708.615 465.119 708.665 465.169 ;
      RECT 708.495 465.119 708.545 465.169 ;
      RECT 708.375 465.119 708.425 465.169 ;
      RECT 708.255 465.119 708.305 465.169 ;
      RECT 708.135 465.119 708.185 465.169 ;
      RECT 708.015 465.119 708.065 465.169 ;
      RECT 707.895 465.119 707.945 465.169 ;
      RECT 707.775 465.119 707.825 465.169 ;
      RECT 707.655 465.119 707.705 465.169 ;
      RECT 707.535 465.119 707.585 465.169 ;
      RECT 646.415 465.119 646.465 465.169 ;
      RECT 646.295 465.119 646.345 465.169 ;
      RECT 646.175 465.119 646.225 465.169 ;
      RECT 646.055 465.119 646.105 465.169 ;
      RECT 645.935 465.119 645.985 465.169 ;
      RECT 645.815 465.119 645.865 465.169 ;
      RECT 645.695 465.119 645.745 465.169 ;
      RECT 645.575 465.119 645.625 465.169 ;
      RECT 645.455 465.119 645.505 465.169 ;
      RECT 645.335 465.119 645.385 465.169 ;
      RECT 645.215 465.119 645.265 465.169 ;
      RECT 645.095 465.119 645.145 465.169 ;
      RECT 644.975 465.119 645.025 465.169 ;
      RECT 644.855 465.119 644.905 465.169 ;
      RECT 644.735 465.119 644.785 465.169 ;
      RECT 644.615 465.119 644.665 465.169 ;
      RECT 644.495 465.119 644.545 465.169 ;
      RECT 644.375 465.119 644.425 465.169 ;
      RECT 644.255 465.119 644.305 465.169 ;
      RECT 644.135 465.119 644.185 465.169 ;
      RECT 644.015 465.119 644.065 465.169 ;
      RECT 643.895 465.119 643.945 465.169 ;
      RECT 643.775 465.119 643.825 465.169 ;
      RECT 643.655 465.119 643.705 465.169 ;
      RECT 643.535 465.119 643.585 465.169 ;
      RECT 576.415 465.119 576.465 465.169 ;
      RECT 576.295 465.119 576.345 465.169 ;
      RECT 576.175 465.119 576.225 465.169 ;
      RECT 576.055 465.119 576.105 465.169 ;
      RECT 575.935 465.119 575.985 465.169 ;
      RECT 575.815 465.119 575.865 465.169 ;
      RECT 575.695 465.119 575.745 465.169 ;
      RECT 575.575 465.119 575.625 465.169 ;
      RECT 575.455 465.119 575.505 465.169 ;
      RECT 575.335 465.119 575.385 465.169 ;
      RECT 575.215 465.119 575.265 465.169 ;
      RECT 575.095 465.119 575.145 465.169 ;
      RECT 574.975 465.119 575.025 465.169 ;
      RECT 574.855 465.119 574.905 465.169 ;
      RECT 574.735 465.119 574.785 465.169 ;
      RECT 574.615 465.119 574.665 465.169 ;
      RECT 574.495 465.119 574.545 465.169 ;
      RECT 574.375 465.119 574.425 465.169 ;
      RECT 574.255 465.119 574.305 465.169 ;
      RECT 574.135 465.119 574.185 465.169 ;
      RECT 574.015 465.119 574.065 465.169 ;
      RECT 573.895 465.119 573.945 465.169 ;
      RECT 573.775 465.119 573.825 465.169 ;
      RECT 573.655 465.119 573.705 465.169 ;
      RECT 573.535 465.119 573.585 465.169 ;
      RECT 510.415 465.119 510.465 465.169 ;
      RECT 510.295 465.119 510.345 465.169 ;
      RECT 510.175 465.119 510.225 465.169 ;
      RECT 510.055 465.119 510.105 465.169 ;
      RECT 509.935 465.119 509.985 465.169 ;
      RECT 509.815 465.119 509.865 465.169 ;
      RECT 509.695 465.119 509.745 465.169 ;
      RECT 509.575 465.119 509.625 465.169 ;
      RECT 509.455 465.119 509.505 465.169 ;
      RECT 509.335 465.119 509.385 465.169 ;
      RECT 509.215 465.119 509.265 465.169 ;
      RECT 509.095 465.119 509.145 465.169 ;
      RECT 508.975 465.119 509.025 465.169 ;
      RECT 508.855 465.119 508.905 465.169 ;
      RECT 508.735 465.119 508.785 465.169 ;
      RECT 508.615 465.119 508.665 465.169 ;
      RECT 508.495 465.119 508.545 465.169 ;
      RECT 508.375 465.119 508.425 465.169 ;
      RECT 508.255 465.119 508.305 465.169 ;
      RECT 508.135 465.119 508.185 465.169 ;
      RECT 508.015 465.119 508.065 465.169 ;
      RECT 507.895 465.119 507.945 465.169 ;
      RECT 507.775 465.119 507.825 465.169 ;
      RECT 507.655 465.119 507.705 465.169 ;
      RECT 507.535 465.119 507.585 465.169 ;
      RECT 446.415 465.119 446.465 465.169 ;
      RECT 446.295 465.119 446.345 465.169 ;
      RECT 446.175 465.119 446.225 465.169 ;
      RECT 446.055 465.119 446.105 465.169 ;
      RECT 445.935 465.119 445.985 465.169 ;
      RECT 445.815 465.119 445.865 465.169 ;
      RECT 445.695 465.119 445.745 465.169 ;
      RECT 445.575 465.119 445.625 465.169 ;
      RECT 445.455 465.119 445.505 465.169 ;
      RECT 445.335 465.119 445.385 465.169 ;
      RECT 445.215 465.119 445.265 465.169 ;
      RECT 445.095 465.119 445.145 465.169 ;
      RECT 444.975 465.119 445.025 465.169 ;
      RECT 444.855 465.119 444.905 465.169 ;
      RECT 444.735 465.119 444.785 465.169 ;
      RECT 444.615 465.119 444.665 465.169 ;
      RECT 444.495 465.119 444.545 465.169 ;
      RECT 444.375 465.119 444.425 465.169 ;
      RECT 444.255 465.119 444.305 465.169 ;
      RECT 444.135 465.119 444.185 465.169 ;
      RECT 444.015 465.119 444.065 465.169 ;
      RECT 443.895 465.119 443.945 465.169 ;
      RECT 443.775 465.119 443.825 465.169 ;
      RECT 443.655 465.119 443.705 465.169 ;
      RECT 443.535 465.119 443.585 465.169 ;
      RECT 376.415 465.119 376.465 465.169 ;
      RECT 376.295 465.119 376.345 465.169 ;
      RECT 376.175 465.119 376.225 465.169 ;
      RECT 376.055 465.119 376.105 465.169 ;
      RECT 375.935 465.119 375.985 465.169 ;
      RECT 375.815 465.119 375.865 465.169 ;
      RECT 375.695 465.119 375.745 465.169 ;
      RECT 375.575 465.119 375.625 465.169 ;
      RECT 375.455 465.119 375.505 465.169 ;
      RECT 375.335 465.119 375.385 465.169 ;
      RECT 375.215 465.119 375.265 465.169 ;
      RECT 375.095 465.119 375.145 465.169 ;
      RECT 374.975 465.119 375.025 465.169 ;
      RECT 374.855 465.119 374.905 465.169 ;
      RECT 374.735 465.119 374.785 465.169 ;
      RECT 374.615 465.119 374.665 465.169 ;
      RECT 374.495 465.119 374.545 465.169 ;
      RECT 374.375 465.119 374.425 465.169 ;
      RECT 374.255 465.119 374.305 465.169 ;
      RECT 374.135 465.119 374.185 465.169 ;
      RECT 374.015 465.119 374.065 465.169 ;
      RECT 373.895 465.119 373.945 465.169 ;
      RECT 373.775 465.119 373.825 465.169 ;
      RECT 373.655 465.119 373.705 465.169 ;
      RECT 373.535 465.119 373.585 465.169 ;
      RECT 310.415 465.119 310.465 465.169 ;
      RECT 310.295 465.119 310.345 465.169 ;
      RECT 310.175 465.119 310.225 465.169 ;
      RECT 310.055 465.119 310.105 465.169 ;
      RECT 309.935 465.119 309.985 465.169 ;
      RECT 309.815 465.119 309.865 465.169 ;
      RECT 309.695 465.119 309.745 465.169 ;
      RECT 309.575 465.119 309.625 465.169 ;
      RECT 309.455 465.119 309.505 465.169 ;
      RECT 309.335 465.119 309.385 465.169 ;
      RECT 309.215 465.119 309.265 465.169 ;
      RECT 309.095 465.119 309.145 465.169 ;
      RECT 308.975 465.119 309.025 465.169 ;
      RECT 308.855 465.119 308.905 465.169 ;
      RECT 308.735 465.119 308.785 465.169 ;
      RECT 308.615 465.119 308.665 465.169 ;
      RECT 308.495 465.119 308.545 465.169 ;
      RECT 308.375 465.119 308.425 465.169 ;
      RECT 308.255 465.119 308.305 465.169 ;
      RECT 308.135 465.119 308.185 465.169 ;
      RECT 308.015 465.119 308.065 465.169 ;
      RECT 307.895 465.119 307.945 465.169 ;
      RECT 307.775 465.119 307.825 465.169 ;
      RECT 307.655 465.119 307.705 465.169 ;
      RECT 307.535 465.119 307.585 465.169 ;
      RECT 246.415 465.119 246.465 465.169 ;
      RECT 246.295 465.119 246.345 465.169 ;
      RECT 246.175 465.119 246.225 465.169 ;
      RECT 246.055 465.119 246.105 465.169 ;
      RECT 245.935 465.119 245.985 465.169 ;
      RECT 245.815 465.119 245.865 465.169 ;
      RECT 245.695 465.119 245.745 465.169 ;
      RECT 245.575 465.119 245.625 465.169 ;
      RECT 245.455 465.119 245.505 465.169 ;
      RECT 245.335 465.119 245.385 465.169 ;
      RECT 245.215 465.119 245.265 465.169 ;
      RECT 245.095 465.119 245.145 465.169 ;
      RECT 244.975 465.119 245.025 465.169 ;
      RECT 244.855 465.119 244.905 465.169 ;
      RECT 244.735 465.119 244.785 465.169 ;
      RECT 244.615 465.119 244.665 465.169 ;
      RECT 244.495 465.119 244.545 465.169 ;
      RECT 244.375 465.119 244.425 465.169 ;
      RECT 244.255 465.119 244.305 465.169 ;
      RECT 244.135 465.119 244.185 465.169 ;
      RECT 244.015 465.119 244.065 465.169 ;
      RECT 243.895 465.119 243.945 465.169 ;
      RECT 243.775 465.119 243.825 465.169 ;
      RECT 243.655 465.119 243.705 465.169 ;
      RECT 243.535 465.119 243.585 465.169 ;
      RECT 176.415 465.119 176.465 465.169 ;
      RECT 176.295 465.119 176.345 465.169 ;
      RECT 176.175 465.119 176.225 465.169 ;
      RECT 176.055 465.119 176.105 465.169 ;
      RECT 175.935 465.119 175.985 465.169 ;
      RECT 175.815 465.119 175.865 465.169 ;
      RECT 175.695 465.119 175.745 465.169 ;
      RECT 175.575 465.119 175.625 465.169 ;
      RECT 175.455 465.119 175.505 465.169 ;
      RECT 175.335 465.119 175.385 465.169 ;
      RECT 175.215 465.119 175.265 465.169 ;
      RECT 175.095 465.119 175.145 465.169 ;
      RECT 174.975 465.119 175.025 465.169 ;
      RECT 174.855 465.119 174.905 465.169 ;
      RECT 174.735 465.119 174.785 465.169 ;
      RECT 174.615 465.119 174.665 465.169 ;
      RECT 174.495 465.119 174.545 465.169 ;
      RECT 174.375 465.119 174.425 465.169 ;
      RECT 174.255 465.119 174.305 465.169 ;
      RECT 174.135 465.119 174.185 465.169 ;
      RECT 174.015 465.119 174.065 465.169 ;
      RECT 173.895 465.119 173.945 465.169 ;
      RECT 173.775 465.119 173.825 465.169 ;
      RECT 173.655 465.119 173.705 465.169 ;
      RECT 173.535 465.119 173.585 465.169 ;
      RECT 110.415 465.119 110.465 465.169 ;
      RECT 110.295 465.119 110.345 465.169 ;
      RECT 110.175 465.119 110.225 465.169 ;
      RECT 110.055 465.119 110.105 465.169 ;
      RECT 109.935 465.119 109.985 465.169 ;
      RECT 109.815 465.119 109.865 465.169 ;
      RECT 109.695 465.119 109.745 465.169 ;
      RECT 109.575 465.119 109.625 465.169 ;
      RECT 109.455 465.119 109.505 465.169 ;
      RECT 109.335 465.119 109.385 465.169 ;
      RECT 109.215 465.119 109.265 465.169 ;
      RECT 109.095 465.119 109.145 465.169 ;
      RECT 108.975 465.119 109.025 465.169 ;
      RECT 108.855 465.119 108.905 465.169 ;
      RECT 108.735 465.119 108.785 465.169 ;
      RECT 108.615 465.119 108.665 465.169 ;
      RECT 108.495 465.119 108.545 465.169 ;
      RECT 108.375 465.119 108.425 465.169 ;
      RECT 108.255 465.119 108.305 465.169 ;
      RECT 108.135 465.119 108.185 465.169 ;
      RECT 108.015 465.119 108.065 465.169 ;
      RECT 107.895 465.119 107.945 465.169 ;
      RECT 107.775 465.119 107.825 465.169 ;
      RECT 107.655 465.119 107.705 465.169 ;
      RECT 107.535 465.119 107.585 465.169 ;
      RECT 46.415 465.119 46.465 465.169 ;
      RECT 46.295 465.119 46.345 465.169 ;
      RECT 46.175 465.119 46.225 465.169 ;
      RECT 46.055 465.119 46.105 465.169 ;
      RECT 45.935 465.119 45.985 465.169 ;
      RECT 45.815 465.119 45.865 465.169 ;
      RECT 45.695 465.119 45.745 465.169 ;
      RECT 45.575 465.119 45.625 465.169 ;
      RECT 45.455 465.119 45.505 465.169 ;
      RECT 45.335 465.119 45.385 465.169 ;
      RECT 45.215 465.119 45.265 465.169 ;
      RECT 45.095 465.119 45.145 465.169 ;
      RECT 44.975 465.119 45.025 465.169 ;
      RECT 44.855 465.119 44.905 465.169 ;
      RECT 44.735 465.119 44.785 465.169 ;
      RECT 44.615 465.119 44.665 465.169 ;
      RECT 44.495 465.119 44.545 465.169 ;
      RECT 44.375 465.119 44.425 465.169 ;
      RECT 44.255 465.119 44.305 465.169 ;
      RECT 44.135 465.119 44.185 465.169 ;
      RECT 44.015 465.119 44.065 465.169 ;
      RECT 43.895 465.119 43.945 465.169 ;
      RECT 43.775 465.119 43.825 465.169 ;
      RECT 43.655 465.119 43.705 465.169 ;
      RECT 43.535 465.119 43.585 465.169 ;
      RECT 1576.415 3.647 1576.465 3.697 ;
      RECT 1576.295 3.647 1576.345 3.697 ;
      RECT 1576.175 3.647 1576.225 3.697 ;
      RECT 1576.055 3.647 1576.105 3.697 ;
      RECT 1575.935 3.647 1575.985 3.697 ;
      RECT 1575.815 3.647 1575.865 3.697 ;
      RECT 1575.695 3.647 1575.745 3.697 ;
      RECT 1575.575 3.647 1575.625 3.697 ;
      RECT 1575.455 3.647 1575.505 3.697 ;
      RECT 1575.335 3.647 1575.385 3.697 ;
      RECT 1575.215 3.647 1575.265 3.697 ;
      RECT 1575.095 3.647 1575.145 3.697 ;
      RECT 1574.975 3.647 1575.025 3.697 ;
      RECT 1574.855 3.647 1574.905 3.697 ;
      RECT 1574.735 3.647 1574.785 3.697 ;
      RECT 1574.615 3.647 1574.665 3.697 ;
      RECT 1574.495 3.647 1574.545 3.697 ;
      RECT 1574.375 3.647 1574.425 3.697 ;
      RECT 1574.255 3.647 1574.305 3.697 ;
      RECT 1574.135 3.647 1574.185 3.697 ;
      RECT 1574.015 3.647 1574.065 3.697 ;
      RECT 1573.895 3.647 1573.945 3.697 ;
      RECT 1573.775 3.647 1573.825 3.697 ;
      RECT 1573.655 3.647 1573.705 3.697 ;
      RECT 1573.535 3.647 1573.585 3.697 ;
      RECT 1510.415 3.647 1510.465 3.697 ;
      RECT 1510.295 3.647 1510.345 3.697 ;
      RECT 1510.175 3.647 1510.225 3.697 ;
      RECT 1510.055 3.647 1510.105 3.697 ;
      RECT 1509.935 3.647 1509.985 3.697 ;
      RECT 1509.815 3.647 1509.865 3.697 ;
      RECT 1509.695 3.647 1509.745 3.697 ;
      RECT 1509.575 3.647 1509.625 3.697 ;
      RECT 1509.455 3.647 1509.505 3.697 ;
      RECT 1509.335 3.647 1509.385 3.697 ;
      RECT 1509.215 3.647 1509.265 3.697 ;
      RECT 1509.095 3.647 1509.145 3.697 ;
      RECT 1508.975 3.647 1509.025 3.697 ;
      RECT 1508.855 3.647 1508.905 3.697 ;
      RECT 1508.735 3.647 1508.785 3.697 ;
      RECT 1508.615 3.647 1508.665 3.697 ;
      RECT 1508.495 3.647 1508.545 3.697 ;
      RECT 1508.375 3.647 1508.425 3.697 ;
      RECT 1508.255 3.647 1508.305 3.697 ;
      RECT 1508.135 3.647 1508.185 3.697 ;
      RECT 1508.015 3.647 1508.065 3.697 ;
      RECT 1507.895 3.647 1507.945 3.697 ;
      RECT 1507.775 3.647 1507.825 3.697 ;
      RECT 1507.655 3.647 1507.705 3.697 ;
      RECT 1507.535 3.647 1507.585 3.697 ;
      RECT 1446.415 3.647 1446.465 3.697 ;
      RECT 1446.295 3.647 1446.345 3.697 ;
      RECT 1446.175 3.647 1446.225 3.697 ;
      RECT 1446.055 3.647 1446.105 3.697 ;
      RECT 1445.935 3.647 1445.985 3.697 ;
      RECT 1445.815 3.647 1445.865 3.697 ;
      RECT 1445.695 3.647 1445.745 3.697 ;
      RECT 1445.575 3.647 1445.625 3.697 ;
      RECT 1445.455 3.647 1445.505 3.697 ;
      RECT 1445.335 3.647 1445.385 3.697 ;
      RECT 1445.215 3.647 1445.265 3.697 ;
      RECT 1445.095 3.647 1445.145 3.697 ;
      RECT 1444.975 3.647 1445.025 3.697 ;
      RECT 1444.855 3.647 1444.905 3.697 ;
      RECT 1444.735 3.647 1444.785 3.697 ;
      RECT 1444.615 3.647 1444.665 3.697 ;
      RECT 1444.495 3.647 1444.545 3.697 ;
      RECT 1444.375 3.647 1444.425 3.697 ;
      RECT 1444.255 3.647 1444.305 3.697 ;
      RECT 1444.135 3.647 1444.185 3.697 ;
      RECT 1444.015 3.647 1444.065 3.697 ;
      RECT 1443.895 3.647 1443.945 3.697 ;
      RECT 1443.775 3.647 1443.825 3.697 ;
      RECT 1443.655 3.647 1443.705 3.697 ;
      RECT 1443.535 3.647 1443.585 3.697 ;
      RECT 1376.415 3.647 1376.465 3.697 ;
      RECT 1376.295 3.647 1376.345 3.697 ;
      RECT 1376.175 3.647 1376.225 3.697 ;
      RECT 1376.055 3.647 1376.105 3.697 ;
      RECT 1375.935 3.647 1375.985 3.697 ;
      RECT 1375.815 3.647 1375.865 3.697 ;
      RECT 1375.695 3.647 1375.745 3.697 ;
      RECT 1375.575 3.647 1375.625 3.697 ;
      RECT 1375.455 3.647 1375.505 3.697 ;
      RECT 1375.335 3.647 1375.385 3.697 ;
      RECT 1375.215 3.647 1375.265 3.697 ;
      RECT 1375.095 3.647 1375.145 3.697 ;
      RECT 1374.975 3.647 1375.025 3.697 ;
      RECT 1374.855 3.647 1374.905 3.697 ;
      RECT 1374.735 3.647 1374.785 3.697 ;
      RECT 1374.615 3.647 1374.665 3.697 ;
      RECT 1374.495 3.647 1374.545 3.697 ;
      RECT 1374.375 3.647 1374.425 3.697 ;
      RECT 1374.255 3.647 1374.305 3.697 ;
      RECT 1374.135 3.647 1374.185 3.697 ;
      RECT 1374.015 3.647 1374.065 3.697 ;
      RECT 1373.895 3.647 1373.945 3.697 ;
      RECT 1373.775 3.647 1373.825 3.697 ;
      RECT 1373.655 3.647 1373.705 3.697 ;
      RECT 1373.535 3.647 1373.585 3.697 ;
      RECT 1310.415 3.647 1310.465 3.697 ;
      RECT 1310.295 3.647 1310.345 3.697 ;
      RECT 1310.175 3.647 1310.225 3.697 ;
      RECT 1310.055 3.647 1310.105 3.697 ;
      RECT 1309.935 3.647 1309.985 3.697 ;
      RECT 1309.815 3.647 1309.865 3.697 ;
      RECT 1309.695 3.647 1309.745 3.697 ;
      RECT 1309.575 3.647 1309.625 3.697 ;
      RECT 1309.455 3.647 1309.505 3.697 ;
      RECT 1309.335 3.647 1309.385 3.697 ;
      RECT 1309.215 3.647 1309.265 3.697 ;
      RECT 1309.095 3.647 1309.145 3.697 ;
      RECT 1308.975 3.647 1309.025 3.697 ;
      RECT 1308.855 3.647 1308.905 3.697 ;
      RECT 1308.735 3.647 1308.785 3.697 ;
      RECT 1308.615 3.647 1308.665 3.697 ;
      RECT 1308.495 3.647 1308.545 3.697 ;
      RECT 1308.375 3.647 1308.425 3.697 ;
      RECT 1308.255 3.647 1308.305 3.697 ;
      RECT 1308.135 3.647 1308.185 3.697 ;
      RECT 1308.015 3.647 1308.065 3.697 ;
      RECT 1307.895 3.647 1307.945 3.697 ;
      RECT 1307.775 3.647 1307.825 3.697 ;
      RECT 1307.655 3.647 1307.705 3.697 ;
      RECT 1307.535 3.647 1307.585 3.697 ;
      RECT 1246.415 3.647 1246.465 3.697 ;
      RECT 1246.295 3.647 1246.345 3.697 ;
      RECT 1246.175 3.647 1246.225 3.697 ;
      RECT 1246.055 3.647 1246.105 3.697 ;
      RECT 1245.935 3.647 1245.985 3.697 ;
      RECT 1245.815 3.647 1245.865 3.697 ;
      RECT 1245.695 3.647 1245.745 3.697 ;
      RECT 1245.575 3.647 1245.625 3.697 ;
      RECT 1245.455 3.647 1245.505 3.697 ;
      RECT 1245.335 3.647 1245.385 3.697 ;
      RECT 1245.215 3.647 1245.265 3.697 ;
      RECT 1245.095 3.647 1245.145 3.697 ;
      RECT 1244.975 3.647 1245.025 3.697 ;
      RECT 1244.855 3.647 1244.905 3.697 ;
      RECT 1244.735 3.647 1244.785 3.697 ;
      RECT 1244.615 3.647 1244.665 3.697 ;
      RECT 1244.495 3.647 1244.545 3.697 ;
      RECT 1244.375 3.647 1244.425 3.697 ;
      RECT 1244.255 3.647 1244.305 3.697 ;
      RECT 1244.135 3.647 1244.185 3.697 ;
      RECT 1244.015 3.647 1244.065 3.697 ;
      RECT 1243.895 3.647 1243.945 3.697 ;
      RECT 1243.775 3.647 1243.825 3.697 ;
      RECT 1243.655 3.647 1243.705 3.697 ;
      RECT 1243.535 3.647 1243.585 3.697 ;
      RECT 1176.415 3.647 1176.465 3.697 ;
      RECT 1176.295 3.647 1176.345 3.697 ;
      RECT 1176.175 3.647 1176.225 3.697 ;
      RECT 1176.055 3.647 1176.105 3.697 ;
      RECT 1175.935 3.647 1175.985 3.697 ;
      RECT 1175.815 3.647 1175.865 3.697 ;
      RECT 1175.695 3.647 1175.745 3.697 ;
      RECT 1175.575 3.647 1175.625 3.697 ;
      RECT 1175.455 3.647 1175.505 3.697 ;
      RECT 1175.335 3.647 1175.385 3.697 ;
      RECT 1175.215 3.647 1175.265 3.697 ;
      RECT 1175.095 3.647 1175.145 3.697 ;
      RECT 1174.975 3.647 1175.025 3.697 ;
      RECT 1174.855 3.647 1174.905 3.697 ;
      RECT 1174.735 3.647 1174.785 3.697 ;
      RECT 1174.615 3.647 1174.665 3.697 ;
      RECT 1174.495 3.647 1174.545 3.697 ;
      RECT 1174.375 3.647 1174.425 3.697 ;
      RECT 1174.255 3.647 1174.305 3.697 ;
      RECT 1174.135 3.647 1174.185 3.697 ;
      RECT 1174.015 3.647 1174.065 3.697 ;
      RECT 1173.895 3.647 1173.945 3.697 ;
      RECT 1173.775 3.647 1173.825 3.697 ;
      RECT 1173.655 3.647 1173.705 3.697 ;
      RECT 1173.535 3.647 1173.585 3.697 ;
      RECT 1110.415 3.647 1110.465 3.697 ;
      RECT 1110.295 3.647 1110.345 3.697 ;
      RECT 1110.175 3.647 1110.225 3.697 ;
      RECT 1110.055 3.647 1110.105 3.697 ;
      RECT 1109.935 3.647 1109.985 3.697 ;
      RECT 1109.815 3.647 1109.865 3.697 ;
      RECT 1109.695 3.647 1109.745 3.697 ;
      RECT 1109.575 3.647 1109.625 3.697 ;
      RECT 1109.455 3.647 1109.505 3.697 ;
      RECT 1109.335 3.647 1109.385 3.697 ;
      RECT 1109.215 3.647 1109.265 3.697 ;
      RECT 1109.095 3.647 1109.145 3.697 ;
      RECT 1108.975 3.647 1109.025 3.697 ;
      RECT 1108.855 3.647 1108.905 3.697 ;
      RECT 1108.735 3.647 1108.785 3.697 ;
      RECT 1108.615 3.647 1108.665 3.697 ;
      RECT 1108.495 3.647 1108.545 3.697 ;
      RECT 1108.375 3.647 1108.425 3.697 ;
      RECT 1108.255 3.647 1108.305 3.697 ;
      RECT 1108.135 3.647 1108.185 3.697 ;
      RECT 1108.015 3.647 1108.065 3.697 ;
      RECT 1107.895 3.647 1107.945 3.697 ;
      RECT 1107.775 3.647 1107.825 3.697 ;
      RECT 1107.655 3.647 1107.705 3.697 ;
      RECT 1107.535 3.647 1107.585 3.697 ;
      RECT 1046.415 3.647 1046.465 3.697 ;
      RECT 1046.295 3.647 1046.345 3.697 ;
      RECT 1046.175 3.647 1046.225 3.697 ;
      RECT 1046.055 3.647 1046.105 3.697 ;
      RECT 1045.935 3.647 1045.985 3.697 ;
      RECT 1045.815 3.647 1045.865 3.697 ;
      RECT 1045.695 3.647 1045.745 3.697 ;
      RECT 1045.575 3.647 1045.625 3.697 ;
      RECT 1045.455 3.647 1045.505 3.697 ;
      RECT 1045.335 3.647 1045.385 3.697 ;
      RECT 1045.215 3.647 1045.265 3.697 ;
      RECT 1045.095 3.647 1045.145 3.697 ;
      RECT 1044.975 3.647 1045.025 3.697 ;
      RECT 1044.855 3.647 1044.905 3.697 ;
      RECT 1044.735 3.647 1044.785 3.697 ;
      RECT 1044.615 3.647 1044.665 3.697 ;
      RECT 1044.495 3.647 1044.545 3.697 ;
      RECT 1044.375 3.647 1044.425 3.697 ;
      RECT 1044.255 3.647 1044.305 3.697 ;
      RECT 1044.135 3.647 1044.185 3.697 ;
      RECT 1044.015 3.647 1044.065 3.697 ;
      RECT 1043.895 3.647 1043.945 3.697 ;
      RECT 1043.775 3.647 1043.825 3.697 ;
      RECT 1043.655 3.647 1043.705 3.697 ;
      RECT 1043.535 3.647 1043.585 3.697 ;
      RECT 976.415 3.647 976.465 3.697 ;
      RECT 976.295 3.647 976.345 3.697 ;
      RECT 976.175 3.647 976.225 3.697 ;
      RECT 976.055 3.647 976.105 3.697 ;
      RECT 975.935 3.647 975.985 3.697 ;
      RECT 975.815 3.647 975.865 3.697 ;
      RECT 975.695 3.647 975.745 3.697 ;
      RECT 975.575 3.647 975.625 3.697 ;
      RECT 975.455 3.647 975.505 3.697 ;
      RECT 975.335 3.647 975.385 3.697 ;
      RECT 975.215 3.647 975.265 3.697 ;
      RECT 975.095 3.647 975.145 3.697 ;
      RECT 974.975 3.647 975.025 3.697 ;
      RECT 974.855 3.647 974.905 3.697 ;
      RECT 974.735 3.647 974.785 3.697 ;
      RECT 974.615 3.647 974.665 3.697 ;
      RECT 974.495 3.647 974.545 3.697 ;
      RECT 974.375 3.647 974.425 3.697 ;
      RECT 974.255 3.647 974.305 3.697 ;
      RECT 974.135 3.647 974.185 3.697 ;
      RECT 974.015 3.647 974.065 3.697 ;
      RECT 973.895 3.647 973.945 3.697 ;
      RECT 973.775 3.647 973.825 3.697 ;
      RECT 973.655 3.647 973.705 3.697 ;
      RECT 973.535 3.647 973.585 3.697 ;
      RECT 910.415 3.647 910.465 3.697 ;
      RECT 910.295 3.647 910.345 3.697 ;
      RECT 910.175 3.647 910.225 3.697 ;
      RECT 910.055 3.647 910.105 3.697 ;
      RECT 909.935 3.647 909.985 3.697 ;
      RECT 909.815 3.647 909.865 3.697 ;
      RECT 909.695 3.647 909.745 3.697 ;
      RECT 909.575 3.647 909.625 3.697 ;
      RECT 909.455 3.647 909.505 3.697 ;
      RECT 909.335 3.647 909.385 3.697 ;
      RECT 909.215 3.647 909.265 3.697 ;
      RECT 909.095 3.647 909.145 3.697 ;
      RECT 908.975 3.647 909.025 3.697 ;
      RECT 908.855 3.647 908.905 3.697 ;
      RECT 908.735 3.647 908.785 3.697 ;
      RECT 908.615 3.647 908.665 3.697 ;
      RECT 908.495 3.647 908.545 3.697 ;
      RECT 908.375 3.647 908.425 3.697 ;
      RECT 908.255 3.647 908.305 3.697 ;
      RECT 908.135 3.647 908.185 3.697 ;
      RECT 908.015 3.647 908.065 3.697 ;
      RECT 907.895 3.647 907.945 3.697 ;
      RECT 907.775 3.647 907.825 3.697 ;
      RECT 907.655 3.647 907.705 3.697 ;
      RECT 907.535 3.647 907.585 3.697 ;
      RECT 846.415 3.647 846.465 3.697 ;
      RECT 846.295 3.647 846.345 3.697 ;
      RECT 846.175 3.647 846.225 3.697 ;
      RECT 846.055 3.647 846.105 3.697 ;
      RECT 845.935 3.647 845.985 3.697 ;
      RECT 845.815 3.647 845.865 3.697 ;
      RECT 845.695 3.647 845.745 3.697 ;
      RECT 845.575 3.647 845.625 3.697 ;
      RECT 845.455 3.647 845.505 3.697 ;
      RECT 845.335 3.647 845.385 3.697 ;
      RECT 845.215 3.647 845.265 3.697 ;
      RECT 845.095 3.647 845.145 3.697 ;
      RECT 844.975 3.647 845.025 3.697 ;
      RECT 844.855 3.647 844.905 3.697 ;
      RECT 844.735 3.647 844.785 3.697 ;
      RECT 844.615 3.647 844.665 3.697 ;
      RECT 844.495 3.647 844.545 3.697 ;
      RECT 844.375 3.647 844.425 3.697 ;
      RECT 844.255 3.647 844.305 3.697 ;
      RECT 844.135 3.647 844.185 3.697 ;
      RECT 844.015 3.647 844.065 3.697 ;
      RECT 843.895 3.647 843.945 3.697 ;
      RECT 843.775 3.647 843.825 3.697 ;
      RECT 843.655 3.647 843.705 3.697 ;
      RECT 843.535 3.647 843.585 3.697 ;
      RECT 776.415 3.647 776.465 3.697 ;
      RECT 776.295 3.647 776.345 3.697 ;
      RECT 776.175 3.647 776.225 3.697 ;
      RECT 776.055 3.647 776.105 3.697 ;
      RECT 775.935 3.647 775.985 3.697 ;
      RECT 775.815 3.647 775.865 3.697 ;
      RECT 775.695 3.647 775.745 3.697 ;
      RECT 775.575 3.647 775.625 3.697 ;
      RECT 775.455 3.647 775.505 3.697 ;
      RECT 775.335 3.647 775.385 3.697 ;
      RECT 775.215 3.647 775.265 3.697 ;
      RECT 775.095 3.647 775.145 3.697 ;
      RECT 774.975 3.647 775.025 3.697 ;
      RECT 774.855 3.647 774.905 3.697 ;
      RECT 774.735 3.647 774.785 3.697 ;
      RECT 774.615 3.647 774.665 3.697 ;
      RECT 774.495 3.647 774.545 3.697 ;
      RECT 774.375 3.647 774.425 3.697 ;
      RECT 774.255 3.647 774.305 3.697 ;
      RECT 774.135 3.647 774.185 3.697 ;
      RECT 774.015 3.647 774.065 3.697 ;
      RECT 773.895 3.647 773.945 3.697 ;
      RECT 773.775 3.647 773.825 3.697 ;
      RECT 773.655 3.647 773.705 3.697 ;
      RECT 773.535 3.647 773.585 3.697 ;
      RECT 710.415 3.647 710.465 3.697 ;
      RECT 710.295 3.647 710.345 3.697 ;
      RECT 710.175 3.647 710.225 3.697 ;
      RECT 710.055 3.647 710.105 3.697 ;
      RECT 709.935 3.647 709.985 3.697 ;
      RECT 709.815 3.647 709.865 3.697 ;
      RECT 709.695 3.647 709.745 3.697 ;
      RECT 709.575 3.647 709.625 3.697 ;
      RECT 709.455 3.647 709.505 3.697 ;
      RECT 709.335 3.647 709.385 3.697 ;
      RECT 709.215 3.647 709.265 3.697 ;
      RECT 709.095 3.647 709.145 3.697 ;
      RECT 708.975 3.647 709.025 3.697 ;
      RECT 708.855 3.647 708.905 3.697 ;
      RECT 708.735 3.647 708.785 3.697 ;
      RECT 708.615 3.647 708.665 3.697 ;
      RECT 708.495 3.647 708.545 3.697 ;
      RECT 708.375 3.647 708.425 3.697 ;
      RECT 708.255 3.647 708.305 3.697 ;
      RECT 708.135 3.647 708.185 3.697 ;
      RECT 708.015 3.647 708.065 3.697 ;
      RECT 707.895 3.647 707.945 3.697 ;
      RECT 707.775 3.647 707.825 3.697 ;
      RECT 707.655 3.647 707.705 3.697 ;
      RECT 707.535 3.647 707.585 3.697 ;
      RECT 646.415 3.647 646.465 3.697 ;
      RECT 646.295 3.647 646.345 3.697 ;
      RECT 646.175 3.647 646.225 3.697 ;
      RECT 646.055 3.647 646.105 3.697 ;
      RECT 645.935 3.647 645.985 3.697 ;
      RECT 645.815 3.647 645.865 3.697 ;
      RECT 645.695 3.647 645.745 3.697 ;
      RECT 645.575 3.647 645.625 3.697 ;
      RECT 645.455 3.647 645.505 3.697 ;
      RECT 645.335 3.647 645.385 3.697 ;
      RECT 645.215 3.647 645.265 3.697 ;
      RECT 645.095 3.647 645.145 3.697 ;
      RECT 644.975 3.647 645.025 3.697 ;
      RECT 644.855 3.647 644.905 3.697 ;
      RECT 644.735 3.647 644.785 3.697 ;
      RECT 644.615 3.647 644.665 3.697 ;
      RECT 644.495 3.647 644.545 3.697 ;
      RECT 644.375 3.647 644.425 3.697 ;
      RECT 644.255 3.647 644.305 3.697 ;
      RECT 644.135 3.647 644.185 3.697 ;
      RECT 644.015 3.647 644.065 3.697 ;
      RECT 643.895 3.647 643.945 3.697 ;
      RECT 643.775 3.647 643.825 3.697 ;
      RECT 643.655 3.647 643.705 3.697 ;
      RECT 643.535 3.647 643.585 3.697 ;
      RECT 576.415 3.647 576.465 3.697 ;
      RECT 576.295 3.647 576.345 3.697 ;
      RECT 576.175 3.647 576.225 3.697 ;
      RECT 576.055 3.647 576.105 3.697 ;
      RECT 575.935 3.647 575.985 3.697 ;
      RECT 575.815 3.647 575.865 3.697 ;
      RECT 575.695 3.647 575.745 3.697 ;
      RECT 575.575 3.647 575.625 3.697 ;
      RECT 575.455 3.647 575.505 3.697 ;
      RECT 575.335 3.647 575.385 3.697 ;
      RECT 575.215 3.647 575.265 3.697 ;
      RECT 575.095 3.647 575.145 3.697 ;
      RECT 574.975 3.647 575.025 3.697 ;
      RECT 574.855 3.647 574.905 3.697 ;
      RECT 574.735 3.647 574.785 3.697 ;
      RECT 574.615 3.647 574.665 3.697 ;
      RECT 574.495 3.647 574.545 3.697 ;
      RECT 574.375 3.647 574.425 3.697 ;
      RECT 574.255 3.647 574.305 3.697 ;
      RECT 574.135 3.647 574.185 3.697 ;
      RECT 574.015 3.647 574.065 3.697 ;
      RECT 573.895 3.647 573.945 3.697 ;
      RECT 573.775 3.647 573.825 3.697 ;
      RECT 573.655 3.647 573.705 3.697 ;
      RECT 573.535 3.647 573.585 3.697 ;
      RECT 510.415 3.647 510.465 3.697 ;
      RECT 510.295 3.647 510.345 3.697 ;
      RECT 510.175 3.647 510.225 3.697 ;
      RECT 510.055 3.647 510.105 3.697 ;
      RECT 509.935 3.647 509.985 3.697 ;
      RECT 509.815 3.647 509.865 3.697 ;
      RECT 509.695 3.647 509.745 3.697 ;
      RECT 509.575 3.647 509.625 3.697 ;
      RECT 509.455 3.647 509.505 3.697 ;
      RECT 509.335 3.647 509.385 3.697 ;
      RECT 509.215 3.647 509.265 3.697 ;
      RECT 509.095 3.647 509.145 3.697 ;
      RECT 508.975 3.647 509.025 3.697 ;
      RECT 508.855 3.647 508.905 3.697 ;
      RECT 508.735 3.647 508.785 3.697 ;
      RECT 508.615 3.647 508.665 3.697 ;
      RECT 508.495 3.647 508.545 3.697 ;
      RECT 508.375 3.647 508.425 3.697 ;
      RECT 508.255 3.647 508.305 3.697 ;
      RECT 508.135 3.647 508.185 3.697 ;
      RECT 508.015 3.647 508.065 3.697 ;
      RECT 507.895 3.647 507.945 3.697 ;
      RECT 507.775 3.647 507.825 3.697 ;
      RECT 507.655 3.647 507.705 3.697 ;
      RECT 507.535 3.647 507.585 3.697 ;
      RECT 446.415 3.647 446.465 3.697 ;
      RECT 446.295 3.647 446.345 3.697 ;
      RECT 446.175 3.647 446.225 3.697 ;
      RECT 446.055 3.647 446.105 3.697 ;
      RECT 445.935 3.647 445.985 3.697 ;
      RECT 445.815 3.647 445.865 3.697 ;
      RECT 445.695 3.647 445.745 3.697 ;
      RECT 445.575 3.647 445.625 3.697 ;
      RECT 445.455 3.647 445.505 3.697 ;
      RECT 445.335 3.647 445.385 3.697 ;
      RECT 445.215 3.647 445.265 3.697 ;
      RECT 445.095 3.647 445.145 3.697 ;
      RECT 444.975 3.647 445.025 3.697 ;
      RECT 444.855 3.647 444.905 3.697 ;
      RECT 444.735 3.647 444.785 3.697 ;
      RECT 444.615 3.647 444.665 3.697 ;
      RECT 444.495 3.647 444.545 3.697 ;
      RECT 444.375 3.647 444.425 3.697 ;
      RECT 444.255 3.647 444.305 3.697 ;
      RECT 444.135 3.647 444.185 3.697 ;
      RECT 444.015 3.647 444.065 3.697 ;
      RECT 443.895 3.647 443.945 3.697 ;
      RECT 443.775 3.647 443.825 3.697 ;
      RECT 443.655 3.647 443.705 3.697 ;
      RECT 443.535 3.647 443.585 3.697 ;
      RECT 376.415 3.647 376.465 3.697 ;
      RECT 376.295 3.647 376.345 3.697 ;
      RECT 376.175 3.647 376.225 3.697 ;
      RECT 376.055 3.647 376.105 3.697 ;
      RECT 375.935 3.647 375.985 3.697 ;
      RECT 375.815 3.647 375.865 3.697 ;
      RECT 375.695 3.647 375.745 3.697 ;
      RECT 375.575 3.647 375.625 3.697 ;
      RECT 375.455 3.647 375.505 3.697 ;
      RECT 375.335 3.647 375.385 3.697 ;
      RECT 375.215 3.647 375.265 3.697 ;
      RECT 375.095 3.647 375.145 3.697 ;
      RECT 374.975 3.647 375.025 3.697 ;
      RECT 374.855 3.647 374.905 3.697 ;
      RECT 374.735 3.647 374.785 3.697 ;
      RECT 374.615 3.647 374.665 3.697 ;
      RECT 374.495 3.647 374.545 3.697 ;
      RECT 374.375 3.647 374.425 3.697 ;
      RECT 374.255 3.647 374.305 3.697 ;
      RECT 374.135 3.647 374.185 3.697 ;
      RECT 374.015 3.647 374.065 3.697 ;
      RECT 373.895 3.647 373.945 3.697 ;
      RECT 373.775 3.647 373.825 3.697 ;
      RECT 373.655 3.647 373.705 3.697 ;
      RECT 373.535 3.647 373.585 3.697 ;
      RECT 310.415 3.647 310.465 3.697 ;
      RECT 310.295 3.647 310.345 3.697 ;
      RECT 310.175 3.647 310.225 3.697 ;
      RECT 310.055 3.647 310.105 3.697 ;
      RECT 309.935 3.647 309.985 3.697 ;
      RECT 309.815 3.647 309.865 3.697 ;
      RECT 309.695 3.647 309.745 3.697 ;
      RECT 309.575 3.647 309.625 3.697 ;
      RECT 309.455 3.647 309.505 3.697 ;
      RECT 309.335 3.647 309.385 3.697 ;
      RECT 309.215 3.647 309.265 3.697 ;
      RECT 309.095 3.647 309.145 3.697 ;
      RECT 308.975 3.647 309.025 3.697 ;
      RECT 308.855 3.647 308.905 3.697 ;
      RECT 308.735 3.647 308.785 3.697 ;
      RECT 308.615 3.647 308.665 3.697 ;
      RECT 308.495 3.647 308.545 3.697 ;
      RECT 308.375 3.647 308.425 3.697 ;
      RECT 308.255 3.647 308.305 3.697 ;
      RECT 308.135 3.647 308.185 3.697 ;
      RECT 308.015 3.647 308.065 3.697 ;
      RECT 307.895 3.647 307.945 3.697 ;
      RECT 307.775 3.647 307.825 3.697 ;
      RECT 307.655 3.647 307.705 3.697 ;
      RECT 307.535 3.647 307.585 3.697 ;
      RECT 246.415 3.647 246.465 3.697 ;
      RECT 246.295 3.647 246.345 3.697 ;
      RECT 246.175 3.647 246.225 3.697 ;
      RECT 246.055 3.647 246.105 3.697 ;
      RECT 245.935 3.647 245.985 3.697 ;
      RECT 245.815 3.647 245.865 3.697 ;
      RECT 245.695 3.647 245.745 3.697 ;
      RECT 245.575 3.647 245.625 3.697 ;
      RECT 245.455 3.647 245.505 3.697 ;
      RECT 245.335 3.647 245.385 3.697 ;
      RECT 245.215 3.647 245.265 3.697 ;
      RECT 245.095 3.647 245.145 3.697 ;
      RECT 244.975 3.647 245.025 3.697 ;
      RECT 244.855 3.647 244.905 3.697 ;
      RECT 244.735 3.647 244.785 3.697 ;
      RECT 244.615 3.647 244.665 3.697 ;
      RECT 244.495 3.647 244.545 3.697 ;
      RECT 244.375 3.647 244.425 3.697 ;
      RECT 244.255 3.647 244.305 3.697 ;
      RECT 244.135 3.647 244.185 3.697 ;
      RECT 244.015 3.647 244.065 3.697 ;
      RECT 243.895 3.647 243.945 3.697 ;
      RECT 243.775 3.647 243.825 3.697 ;
      RECT 243.655 3.647 243.705 3.697 ;
      RECT 243.535 3.647 243.585 3.697 ;
      RECT 176.415 3.647 176.465 3.697 ;
      RECT 176.295 3.647 176.345 3.697 ;
      RECT 176.175 3.647 176.225 3.697 ;
      RECT 176.055 3.647 176.105 3.697 ;
      RECT 175.935 3.647 175.985 3.697 ;
      RECT 175.815 3.647 175.865 3.697 ;
      RECT 175.695 3.647 175.745 3.697 ;
      RECT 175.575 3.647 175.625 3.697 ;
      RECT 175.455 3.647 175.505 3.697 ;
      RECT 175.335 3.647 175.385 3.697 ;
      RECT 175.215 3.647 175.265 3.697 ;
      RECT 175.095 3.647 175.145 3.697 ;
      RECT 174.975 3.647 175.025 3.697 ;
      RECT 174.855 3.647 174.905 3.697 ;
      RECT 174.735 3.647 174.785 3.697 ;
      RECT 174.615 3.647 174.665 3.697 ;
      RECT 174.495 3.647 174.545 3.697 ;
      RECT 174.375 3.647 174.425 3.697 ;
      RECT 174.255 3.647 174.305 3.697 ;
      RECT 174.135 3.647 174.185 3.697 ;
      RECT 174.015 3.647 174.065 3.697 ;
      RECT 173.895 3.647 173.945 3.697 ;
      RECT 173.775 3.647 173.825 3.697 ;
      RECT 173.655 3.647 173.705 3.697 ;
      RECT 173.535 3.647 173.585 3.697 ;
      RECT 110.415 3.647 110.465 3.697 ;
      RECT 110.295 3.647 110.345 3.697 ;
      RECT 110.175 3.647 110.225 3.697 ;
      RECT 110.055 3.647 110.105 3.697 ;
      RECT 109.935 3.647 109.985 3.697 ;
      RECT 109.815 3.647 109.865 3.697 ;
      RECT 109.695 3.647 109.745 3.697 ;
      RECT 109.575 3.647 109.625 3.697 ;
      RECT 109.455 3.647 109.505 3.697 ;
      RECT 109.335 3.647 109.385 3.697 ;
      RECT 109.215 3.647 109.265 3.697 ;
      RECT 109.095 3.647 109.145 3.697 ;
      RECT 108.975 3.647 109.025 3.697 ;
      RECT 108.855 3.647 108.905 3.697 ;
      RECT 108.735 3.647 108.785 3.697 ;
      RECT 108.615 3.647 108.665 3.697 ;
      RECT 108.495 3.647 108.545 3.697 ;
      RECT 108.375 3.647 108.425 3.697 ;
      RECT 108.255 3.647 108.305 3.697 ;
      RECT 108.135 3.647 108.185 3.697 ;
      RECT 108.015 3.647 108.065 3.697 ;
      RECT 107.895 3.647 107.945 3.697 ;
      RECT 107.775 3.647 107.825 3.697 ;
      RECT 107.655 3.647 107.705 3.697 ;
      RECT 107.535 3.647 107.585 3.697 ;
      RECT 46.415 3.647 46.465 3.697 ;
      RECT 46.295 3.647 46.345 3.697 ;
      RECT 46.175 3.647 46.225 3.697 ;
      RECT 46.055 3.647 46.105 3.697 ;
      RECT 45.935 3.647 45.985 3.697 ;
      RECT 45.815 3.647 45.865 3.697 ;
      RECT 45.695 3.647 45.745 3.697 ;
      RECT 45.575 3.647 45.625 3.697 ;
      RECT 45.455 3.647 45.505 3.697 ;
      RECT 45.335 3.647 45.385 3.697 ;
      RECT 45.215 3.647 45.265 3.697 ;
      RECT 45.095 3.647 45.145 3.697 ;
      RECT 44.975 3.647 45.025 3.697 ;
      RECT 44.855 3.647 44.905 3.697 ;
      RECT 44.735 3.647 44.785 3.697 ;
      RECT 44.615 3.647 44.665 3.697 ;
      RECT 44.495 3.647 44.545 3.697 ;
      RECT 44.375 3.647 44.425 3.697 ;
      RECT 44.255 3.647 44.305 3.697 ;
      RECT 44.135 3.647 44.185 3.697 ;
      RECT 44.015 3.647 44.065 3.697 ;
      RECT 43.895 3.647 43.945 3.697 ;
      RECT 43.775 3.647 43.825 3.697 ;
      RECT 43.655 3.647 43.705 3.697 ;
      RECT 43.535 3.647 43.585 3.697 ;
      RECT 1571.415 1.975 1571.465 2.025 ;
      RECT 1571.295 1.975 1571.345 2.025 ;
      RECT 1571.175 1.975 1571.225 2.025 ;
      RECT 1571.055 1.975 1571.105 2.025 ;
      RECT 1570.935 1.975 1570.985 2.025 ;
      RECT 1570.815 1.975 1570.865 2.025 ;
      RECT 1570.695 1.975 1570.745 2.025 ;
      RECT 1570.575 1.975 1570.625 2.025 ;
      RECT 1570.455 1.975 1570.505 2.025 ;
      RECT 1570.335 1.975 1570.385 2.025 ;
      RECT 1570.215 1.975 1570.265 2.025 ;
      RECT 1570.095 1.975 1570.145 2.025 ;
      RECT 1569.975 1.975 1570.025 2.025 ;
      RECT 1569.855 1.975 1569.905 2.025 ;
      RECT 1569.735 1.975 1569.785 2.025 ;
      RECT 1569.615 1.975 1569.665 2.025 ;
      RECT 1569.495 1.975 1569.545 2.025 ;
      RECT 1569.375 1.975 1569.425 2.025 ;
      RECT 1569.255 1.975 1569.305 2.025 ;
      RECT 1569.135 1.975 1569.185 2.025 ;
      RECT 1569.015 1.975 1569.065 2.025 ;
      RECT 1568.895 1.975 1568.945 2.025 ;
      RECT 1568.775 1.975 1568.825 2.025 ;
      RECT 1568.655 1.975 1568.705 2.025 ;
      RECT 1568.535 1.975 1568.585 2.025 ;
      RECT 1505.415 1.975 1505.465 2.025 ;
      RECT 1505.295 1.975 1505.345 2.025 ;
      RECT 1505.175 1.975 1505.225 2.025 ;
      RECT 1505.055 1.975 1505.105 2.025 ;
      RECT 1504.935 1.975 1504.985 2.025 ;
      RECT 1504.815 1.975 1504.865 2.025 ;
      RECT 1504.695 1.975 1504.745 2.025 ;
      RECT 1504.575 1.975 1504.625 2.025 ;
      RECT 1504.455 1.975 1504.505 2.025 ;
      RECT 1504.335 1.975 1504.385 2.025 ;
      RECT 1504.215 1.975 1504.265 2.025 ;
      RECT 1504.095 1.975 1504.145 2.025 ;
      RECT 1503.975 1.975 1504.025 2.025 ;
      RECT 1503.855 1.975 1503.905 2.025 ;
      RECT 1503.735 1.975 1503.785 2.025 ;
      RECT 1503.615 1.975 1503.665 2.025 ;
      RECT 1503.495 1.975 1503.545 2.025 ;
      RECT 1503.375 1.975 1503.425 2.025 ;
      RECT 1503.255 1.975 1503.305 2.025 ;
      RECT 1503.135 1.975 1503.185 2.025 ;
      RECT 1503.015 1.975 1503.065 2.025 ;
      RECT 1502.895 1.975 1502.945 2.025 ;
      RECT 1502.775 1.975 1502.825 2.025 ;
      RECT 1502.655 1.975 1502.705 2.025 ;
      RECT 1502.535 1.975 1502.585 2.025 ;
      RECT 1441.415 1.975 1441.465 2.025 ;
      RECT 1441.295 1.975 1441.345 2.025 ;
      RECT 1441.175 1.975 1441.225 2.025 ;
      RECT 1441.055 1.975 1441.105 2.025 ;
      RECT 1440.935 1.975 1440.985 2.025 ;
      RECT 1440.815 1.975 1440.865 2.025 ;
      RECT 1440.695 1.975 1440.745 2.025 ;
      RECT 1440.575 1.975 1440.625 2.025 ;
      RECT 1440.455 1.975 1440.505 2.025 ;
      RECT 1440.335 1.975 1440.385 2.025 ;
      RECT 1440.215 1.975 1440.265 2.025 ;
      RECT 1440.095 1.975 1440.145 2.025 ;
      RECT 1439.975 1.975 1440.025 2.025 ;
      RECT 1439.855 1.975 1439.905 2.025 ;
      RECT 1439.735 1.975 1439.785 2.025 ;
      RECT 1439.615 1.975 1439.665 2.025 ;
      RECT 1439.495 1.975 1439.545 2.025 ;
      RECT 1439.375 1.975 1439.425 2.025 ;
      RECT 1439.255 1.975 1439.305 2.025 ;
      RECT 1439.135 1.975 1439.185 2.025 ;
      RECT 1439.015 1.975 1439.065 2.025 ;
      RECT 1438.895 1.975 1438.945 2.025 ;
      RECT 1438.775 1.975 1438.825 2.025 ;
      RECT 1438.655 1.975 1438.705 2.025 ;
      RECT 1438.535 1.975 1438.585 2.025 ;
      RECT 1371.415 1.975 1371.465 2.025 ;
      RECT 1371.295 1.975 1371.345 2.025 ;
      RECT 1371.175 1.975 1371.225 2.025 ;
      RECT 1371.055 1.975 1371.105 2.025 ;
      RECT 1370.935 1.975 1370.985 2.025 ;
      RECT 1370.815 1.975 1370.865 2.025 ;
      RECT 1370.695 1.975 1370.745 2.025 ;
      RECT 1370.575 1.975 1370.625 2.025 ;
      RECT 1370.455 1.975 1370.505 2.025 ;
      RECT 1370.335 1.975 1370.385 2.025 ;
      RECT 1370.215 1.975 1370.265 2.025 ;
      RECT 1370.095 1.975 1370.145 2.025 ;
      RECT 1369.975 1.975 1370.025 2.025 ;
      RECT 1369.855 1.975 1369.905 2.025 ;
      RECT 1369.735 1.975 1369.785 2.025 ;
      RECT 1369.615 1.975 1369.665 2.025 ;
      RECT 1369.495 1.975 1369.545 2.025 ;
      RECT 1369.375 1.975 1369.425 2.025 ;
      RECT 1369.255 1.975 1369.305 2.025 ;
      RECT 1369.135 1.975 1369.185 2.025 ;
      RECT 1369.015 1.975 1369.065 2.025 ;
      RECT 1368.895 1.975 1368.945 2.025 ;
      RECT 1368.775 1.975 1368.825 2.025 ;
      RECT 1368.655 1.975 1368.705 2.025 ;
      RECT 1368.535 1.975 1368.585 2.025 ;
      RECT 1305.415 1.975 1305.465 2.025 ;
      RECT 1305.295 1.975 1305.345 2.025 ;
      RECT 1305.175 1.975 1305.225 2.025 ;
      RECT 1305.055 1.975 1305.105 2.025 ;
      RECT 1304.935 1.975 1304.985 2.025 ;
      RECT 1304.815 1.975 1304.865 2.025 ;
      RECT 1304.695 1.975 1304.745 2.025 ;
      RECT 1304.575 1.975 1304.625 2.025 ;
      RECT 1304.455 1.975 1304.505 2.025 ;
      RECT 1304.335 1.975 1304.385 2.025 ;
      RECT 1304.215 1.975 1304.265 2.025 ;
      RECT 1304.095 1.975 1304.145 2.025 ;
      RECT 1303.975 1.975 1304.025 2.025 ;
      RECT 1303.855 1.975 1303.905 2.025 ;
      RECT 1303.735 1.975 1303.785 2.025 ;
      RECT 1303.615 1.975 1303.665 2.025 ;
      RECT 1303.495 1.975 1303.545 2.025 ;
      RECT 1303.375 1.975 1303.425 2.025 ;
      RECT 1303.255 1.975 1303.305 2.025 ;
      RECT 1303.135 1.975 1303.185 2.025 ;
      RECT 1303.015 1.975 1303.065 2.025 ;
      RECT 1302.895 1.975 1302.945 2.025 ;
      RECT 1302.775 1.975 1302.825 2.025 ;
      RECT 1302.655 1.975 1302.705 2.025 ;
      RECT 1302.535 1.975 1302.585 2.025 ;
      RECT 1241.415 1.975 1241.465 2.025 ;
      RECT 1241.295 1.975 1241.345 2.025 ;
      RECT 1241.175 1.975 1241.225 2.025 ;
      RECT 1241.055 1.975 1241.105 2.025 ;
      RECT 1240.935 1.975 1240.985 2.025 ;
      RECT 1240.815 1.975 1240.865 2.025 ;
      RECT 1240.695 1.975 1240.745 2.025 ;
      RECT 1240.575 1.975 1240.625 2.025 ;
      RECT 1240.455 1.975 1240.505 2.025 ;
      RECT 1240.335 1.975 1240.385 2.025 ;
      RECT 1240.215 1.975 1240.265 2.025 ;
      RECT 1240.095 1.975 1240.145 2.025 ;
      RECT 1239.975 1.975 1240.025 2.025 ;
      RECT 1239.855 1.975 1239.905 2.025 ;
      RECT 1239.735 1.975 1239.785 2.025 ;
      RECT 1239.615 1.975 1239.665 2.025 ;
      RECT 1239.495 1.975 1239.545 2.025 ;
      RECT 1239.375 1.975 1239.425 2.025 ;
      RECT 1239.255 1.975 1239.305 2.025 ;
      RECT 1239.135 1.975 1239.185 2.025 ;
      RECT 1239.015 1.975 1239.065 2.025 ;
      RECT 1238.895 1.975 1238.945 2.025 ;
      RECT 1238.775 1.975 1238.825 2.025 ;
      RECT 1238.655 1.975 1238.705 2.025 ;
      RECT 1238.535 1.975 1238.585 2.025 ;
      RECT 1171.415 1.975 1171.465 2.025 ;
      RECT 1171.295 1.975 1171.345 2.025 ;
      RECT 1171.175 1.975 1171.225 2.025 ;
      RECT 1171.055 1.975 1171.105 2.025 ;
      RECT 1170.935 1.975 1170.985 2.025 ;
      RECT 1170.815 1.975 1170.865 2.025 ;
      RECT 1170.695 1.975 1170.745 2.025 ;
      RECT 1170.575 1.975 1170.625 2.025 ;
      RECT 1170.455 1.975 1170.505 2.025 ;
      RECT 1170.335 1.975 1170.385 2.025 ;
      RECT 1170.215 1.975 1170.265 2.025 ;
      RECT 1170.095 1.975 1170.145 2.025 ;
      RECT 1169.975 1.975 1170.025 2.025 ;
      RECT 1169.855 1.975 1169.905 2.025 ;
      RECT 1169.735 1.975 1169.785 2.025 ;
      RECT 1169.615 1.975 1169.665 2.025 ;
      RECT 1169.495 1.975 1169.545 2.025 ;
      RECT 1169.375 1.975 1169.425 2.025 ;
      RECT 1169.255 1.975 1169.305 2.025 ;
      RECT 1169.135 1.975 1169.185 2.025 ;
      RECT 1169.015 1.975 1169.065 2.025 ;
      RECT 1168.895 1.975 1168.945 2.025 ;
      RECT 1168.775 1.975 1168.825 2.025 ;
      RECT 1168.655 1.975 1168.705 2.025 ;
      RECT 1168.535 1.975 1168.585 2.025 ;
      RECT 1105.415 1.975 1105.465 2.025 ;
      RECT 1105.295 1.975 1105.345 2.025 ;
      RECT 1105.175 1.975 1105.225 2.025 ;
      RECT 1105.055 1.975 1105.105 2.025 ;
      RECT 1104.935 1.975 1104.985 2.025 ;
      RECT 1104.815 1.975 1104.865 2.025 ;
      RECT 1104.695 1.975 1104.745 2.025 ;
      RECT 1104.575 1.975 1104.625 2.025 ;
      RECT 1104.455 1.975 1104.505 2.025 ;
      RECT 1104.335 1.975 1104.385 2.025 ;
      RECT 1104.215 1.975 1104.265 2.025 ;
      RECT 1104.095 1.975 1104.145 2.025 ;
      RECT 1103.975 1.975 1104.025 2.025 ;
      RECT 1103.855 1.975 1103.905 2.025 ;
      RECT 1103.735 1.975 1103.785 2.025 ;
      RECT 1103.615 1.975 1103.665 2.025 ;
      RECT 1103.495 1.975 1103.545 2.025 ;
      RECT 1103.375 1.975 1103.425 2.025 ;
      RECT 1103.255 1.975 1103.305 2.025 ;
      RECT 1103.135 1.975 1103.185 2.025 ;
      RECT 1103.015 1.975 1103.065 2.025 ;
      RECT 1102.895 1.975 1102.945 2.025 ;
      RECT 1102.775 1.975 1102.825 2.025 ;
      RECT 1102.655 1.975 1102.705 2.025 ;
      RECT 1102.535 1.975 1102.585 2.025 ;
      RECT 1041.415 1.975 1041.465 2.025 ;
      RECT 1041.295 1.975 1041.345 2.025 ;
      RECT 1041.175 1.975 1041.225 2.025 ;
      RECT 1041.055 1.975 1041.105 2.025 ;
      RECT 1040.935 1.975 1040.985 2.025 ;
      RECT 1040.815 1.975 1040.865 2.025 ;
      RECT 1040.695 1.975 1040.745 2.025 ;
      RECT 1040.575 1.975 1040.625 2.025 ;
      RECT 1040.455 1.975 1040.505 2.025 ;
      RECT 1040.335 1.975 1040.385 2.025 ;
      RECT 1040.215 1.975 1040.265 2.025 ;
      RECT 1040.095 1.975 1040.145 2.025 ;
      RECT 1039.975 1.975 1040.025 2.025 ;
      RECT 1039.855 1.975 1039.905 2.025 ;
      RECT 1039.735 1.975 1039.785 2.025 ;
      RECT 1039.615 1.975 1039.665 2.025 ;
      RECT 1039.495 1.975 1039.545 2.025 ;
      RECT 1039.375 1.975 1039.425 2.025 ;
      RECT 1039.255 1.975 1039.305 2.025 ;
      RECT 1039.135 1.975 1039.185 2.025 ;
      RECT 1039.015 1.975 1039.065 2.025 ;
      RECT 1038.895 1.975 1038.945 2.025 ;
      RECT 1038.775 1.975 1038.825 2.025 ;
      RECT 1038.655 1.975 1038.705 2.025 ;
      RECT 1038.535 1.975 1038.585 2.025 ;
      RECT 971.415 1.975 971.465 2.025 ;
      RECT 971.295 1.975 971.345 2.025 ;
      RECT 971.175 1.975 971.225 2.025 ;
      RECT 971.055 1.975 971.105 2.025 ;
      RECT 970.935 1.975 970.985 2.025 ;
      RECT 970.815 1.975 970.865 2.025 ;
      RECT 970.695 1.975 970.745 2.025 ;
      RECT 970.575 1.975 970.625 2.025 ;
      RECT 970.455 1.975 970.505 2.025 ;
      RECT 970.335 1.975 970.385 2.025 ;
      RECT 970.215 1.975 970.265 2.025 ;
      RECT 970.095 1.975 970.145 2.025 ;
      RECT 969.975 1.975 970.025 2.025 ;
      RECT 969.855 1.975 969.905 2.025 ;
      RECT 969.735 1.975 969.785 2.025 ;
      RECT 969.615 1.975 969.665 2.025 ;
      RECT 969.495 1.975 969.545 2.025 ;
      RECT 969.375 1.975 969.425 2.025 ;
      RECT 969.255 1.975 969.305 2.025 ;
      RECT 969.135 1.975 969.185 2.025 ;
      RECT 969.015 1.975 969.065 2.025 ;
      RECT 968.895 1.975 968.945 2.025 ;
      RECT 968.775 1.975 968.825 2.025 ;
      RECT 968.655 1.975 968.705 2.025 ;
      RECT 968.535 1.975 968.585 2.025 ;
      RECT 905.415 1.975 905.465 2.025 ;
      RECT 905.295 1.975 905.345 2.025 ;
      RECT 905.175 1.975 905.225 2.025 ;
      RECT 905.055 1.975 905.105 2.025 ;
      RECT 904.935 1.975 904.985 2.025 ;
      RECT 904.815 1.975 904.865 2.025 ;
      RECT 904.695 1.975 904.745 2.025 ;
      RECT 904.575 1.975 904.625 2.025 ;
      RECT 904.455 1.975 904.505 2.025 ;
      RECT 904.335 1.975 904.385 2.025 ;
      RECT 904.215 1.975 904.265 2.025 ;
      RECT 904.095 1.975 904.145 2.025 ;
      RECT 903.975 1.975 904.025 2.025 ;
      RECT 903.855 1.975 903.905 2.025 ;
      RECT 903.735 1.975 903.785 2.025 ;
      RECT 903.615 1.975 903.665 2.025 ;
      RECT 903.495 1.975 903.545 2.025 ;
      RECT 903.375 1.975 903.425 2.025 ;
      RECT 903.255 1.975 903.305 2.025 ;
      RECT 903.135 1.975 903.185 2.025 ;
      RECT 903.015 1.975 903.065 2.025 ;
      RECT 902.895 1.975 902.945 2.025 ;
      RECT 902.775 1.975 902.825 2.025 ;
      RECT 902.655 1.975 902.705 2.025 ;
      RECT 902.535 1.975 902.585 2.025 ;
      RECT 841.415 1.975 841.465 2.025 ;
      RECT 841.295 1.975 841.345 2.025 ;
      RECT 841.175 1.975 841.225 2.025 ;
      RECT 841.055 1.975 841.105 2.025 ;
      RECT 840.935 1.975 840.985 2.025 ;
      RECT 840.815 1.975 840.865 2.025 ;
      RECT 840.695 1.975 840.745 2.025 ;
      RECT 840.575 1.975 840.625 2.025 ;
      RECT 840.455 1.975 840.505 2.025 ;
      RECT 840.335 1.975 840.385 2.025 ;
      RECT 840.215 1.975 840.265 2.025 ;
      RECT 840.095 1.975 840.145 2.025 ;
      RECT 839.975 1.975 840.025 2.025 ;
      RECT 839.855 1.975 839.905 2.025 ;
      RECT 839.735 1.975 839.785 2.025 ;
      RECT 839.615 1.975 839.665 2.025 ;
      RECT 839.495 1.975 839.545 2.025 ;
      RECT 839.375 1.975 839.425 2.025 ;
      RECT 839.255 1.975 839.305 2.025 ;
      RECT 839.135 1.975 839.185 2.025 ;
      RECT 839.015 1.975 839.065 2.025 ;
      RECT 838.895 1.975 838.945 2.025 ;
      RECT 838.775 1.975 838.825 2.025 ;
      RECT 838.655 1.975 838.705 2.025 ;
      RECT 838.535 1.975 838.585 2.025 ;
      RECT 771.415 1.975 771.465 2.025 ;
      RECT 771.295 1.975 771.345 2.025 ;
      RECT 771.175 1.975 771.225 2.025 ;
      RECT 771.055 1.975 771.105 2.025 ;
      RECT 770.935 1.975 770.985 2.025 ;
      RECT 770.815 1.975 770.865 2.025 ;
      RECT 770.695 1.975 770.745 2.025 ;
      RECT 770.575 1.975 770.625 2.025 ;
      RECT 770.455 1.975 770.505 2.025 ;
      RECT 770.335 1.975 770.385 2.025 ;
      RECT 770.215 1.975 770.265 2.025 ;
      RECT 770.095 1.975 770.145 2.025 ;
      RECT 769.975 1.975 770.025 2.025 ;
      RECT 769.855 1.975 769.905 2.025 ;
      RECT 769.735 1.975 769.785 2.025 ;
      RECT 769.615 1.975 769.665 2.025 ;
      RECT 769.495 1.975 769.545 2.025 ;
      RECT 769.375 1.975 769.425 2.025 ;
      RECT 769.255 1.975 769.305 2.025 ;
      RECT 769.135 1.975 769.185 2.025 ;
      RECT 769.015 1.975 769.065 2.025 ;
      RECT 768.895 1.975 768.945 2.025 ;
      RECT 768.775 1.975 768.825 2.025 ;
      RECT 768.655 1.975 768.705 2.025 ;
      RECT 768.535 1.975 768.585 2.025 ;
      RECT 705.415 1.975 705.465 2.025 ;
      RECT 705.295 1.975 705.345 2.025 ;
      RECT 705.175 1.975 705.225 2.025 ;
      RECT 705.055 1.975 705.105 2.025 ;
      RECT 704.935 1.975 704.985 2.025 ;
      RECT 704.815 1.975 704.865 2.025 ;
      RECT 704.695 1.975 704.745 2.025 ;
      RECT 704.575 1.975 704.625 2.025 ;
      RECT 704.455 1.975 704.505 2.025 ;
      RECT 704.335 1.975 704.385 2.025 ;
      RECT 704.215 1.975 704.265 2.025 ;
      RECT 704.095 1.975 704.145 2.025 ;
      RECT 703.975 1.975 704.025 2.025 ;
      RECT 703.855 1.975 703.905 2.025 ;
      RECT 703.735 1.975 703.785 2.025 ;
      RECT 703.615 1.975 703.665 2.025 ;
      RECT 703.495 1.975 703.545 2.025 ;
      RECT 703.375 1.975 703.425 2.025 ;
      RECT 703.255 1.975 703.305 2.025 ;
      RECT 703.135 1.975 703.185 2.025 ;
      RECT 703.015 1.975 703.065 2.025 ;
      RECT 702.895 1.975 702.945 2.025 ;
      RECT 702.775 1.975 702.825 2.025 ;
      RECT 702.655 1.975 702.705 2.025 ;
      RECT 702.535 1.975 702.585 2.025 ;
      RECT 641.415 1.975 641.465 2.025 ;
      RECT 641.295 1.975 641.345 2.025 ;
      RECT 641.175 1.975 641.225 2.025 ;
      RECT 641.055 1.975 641.105 2.025 ;
      RECT 640.935 1.975 640.985 2.025 ;
      RECT 640.815 1.975 640.865 2.025 ;
      RECT 640.695 1.975 640.745 2.025 ;
      RECT 640.575 1.975 640.625 2.025 ;
      RECT 640.455 1.975 640.505 2.025 ;
      RECT 640.335 1.975 640.385 2.025 ;
      RECT 640.215 1.975 640.265 2.025 ;
      RECT 640.095 1.975 640.145 2.025 ;
      RECT 639.975 1.975 640.025 2.025 ;
      RECT 639.855 1.975 639.905 2.025 ;
      RECT 639.735 1.975 639.785 2.025 ;
      RECT 639.615 1.975 639.665 2.025 ;
      RECT 639.495 1.975 639.545 2.025 ;
      RECT 639.375 1.975 639.425 2.025 ;
      RECT 639.255 1.975 639.305 2.025 ;
      RECT 639.135 1.975 639.185 2.025 ;
      RECT 639.015 1.975 639.065 2.025 ;
      RECT 638.895 1.975 638.945 2.025 ;
      RECT 638.775 1.975 638.825 2.025 ;
      RECT 638.655 1.975 638.705 2.025 ;
      RECT 638.535 1.975 638.585 2.025 ;
      RECT 571.415 1.975 571.465 2.025 ;
      RECT 571.295 1.975 571.345 2.025 ;
      RECT 571.175 1.975 571.225 2.025 ;
      RECT 571.055 1.975 571.105 2.025 ;
      RECT 570.935 1.975 570.985 2.025 ;
      RECT 570.815 1.975 570.865 2.025 ;
      RECT 570.695 1.975 570.745 2.025 ;
      RECT 570.575 1.975 570.625 2.025 ;
      RECT 570.455 1.975 570.505 2.025 ;
      RECT 570.335 1.975 570.385 2.025 ;
      RECT 570.215 1.975 570.265 2.025 ;
      RECT 570.095 1.975 570.145 2.025 ;
      RECT 569.975 1.975 570.025 2.025 ;
      RECT 569.855 1.975 569.905 2.025 ;
      RECT 569.735 1.975 569.785 2.025 ;
      RECT 569.615 1.975 569.665 2.025 ;
      RECT 569.495 1.975 569.545 2.025 ;
      RECT 569.375 1.975 569.425 2.025 ;
      RECT 569.255 1.975 569.305 2.025 ;
      RECT 569.135 1.975 569.185 2.025 ;
      RECT 569.015 1.975 569.065 2.025 ;
      RECT 568.895 1.975 568.945 2.025 ;
      RECT 568.775 1.975 568.825 2.025 ;
      RECT 568.655 1.975 568.705 2.025 ;
      RECT 568.535 1.975 568.585 2.025 ;
      RECT 505.415 1.975 505.465 2.025 ;
      RECT 505.295 1.975 505.345 2.025 ;
      RECT 505.175 1.975 505.225 2.025 ;
      RECT 505.055 1.975 505.105 2.025 ;
      RECT 504.935 1.975 504.985 2.025 ;
      RECT 504.815 1.975 504.865 2.025 ;
      RECT 504.695 1.975 504.745 2.025 ;
      RECT 504.575 1.975 504.625 2.025 ;
      RECT 504.455 1.975 504.505 2.025 ;
      RECT 504.335 1.975 504.385 2.025 ;
      RECT 504.215 1.975 504.265 2.025 ;
      RECT 504.095 1.975 504.145 2.025 ;
      RECT 503.975 1.975 504.025 2.025 ;
      RECT 503.855 1.975 503.905 2.025 ;
      RECT 503.735 1.975 503.785 2.025 ;
      RECT 503.615 1.975 503.665 2.025 ;
      RECT 503.495 1.975 503.545 2.025 ;
      RECT 503.375 1.975 503.425 2.025 ;
      RECT 503.255 1.975 503.305 2.025 ;
      RECT 503.135 1.975 503.185 2.025 ;
      RECT 503.015 1.975 503.065 2.025 ;
      RECT 502.895 1.975 502.945 2.025 ;
      RECT 502.775 1.975 502.825 2.025 ;
      RECT 502.655 1.975 502.705 2.025 ;
      RECT 502.535 1.975 502.585 2.025 ;
      RECT 441.415 1.975 441.465 2.025 ;
      RECT 441.295 1.975 441.345 2.025 ;
      RECT 441.175 1.975 441.225 2.025 ;
      RECT 441.055 1.975 441.105 2.025 ;
      RECT 440.935 1.975 440.985 2.025 ;
      RECT 440.815 1.975 440.865 2.025 ;
      RECT 440.695 1.975 440.745 2.025 ;
      RECT 440.575 1.975 440.625 2.025 ;
      RECT 440.455 1.975 440.505 2.025 ;
      RECT 440.335 1.975 440.385 2.025 ;
      RECT 440.215 1.975 440.265 2.025 ;
      RECT 440.095 1.975 440.145 2.025 ;
      RECT 439.975 1.975 440.025 2.025 ;
      RECT 439.855 1.975 439.905 2.025 ;
      RECT 439.735 1.975 439.785 2.025 ;
      RECT 439.615 1.975 439.665 2.025 ;
      RECT 439.495 1.975 439.545 2.025 ;
      RECT 439.375 1.975 439.425 2.025 ;
      RECT 439.255 1.975 439.305 2.025 ;
      RECT 439.135 1.975 439.185 2.025 ;
      RECT 439.015 1.975 439.065 2.025 ;
      RECT 438.895 1.975 438.945 2.025 ;
      RECT 438.775 1.975 438.825 2.025 ;
      RECT 438.655 1.975 438.705 2.025 ;
      RECT 438.535 1.975 438.585 2.025 ;
      RECT 371.415 1.975 371.465 2.025 ;
      RECT 371.295 1.975 371.345 2.025 ;
      RECT 371.175 1.975 371.225 2.025 ;
      RECT 371.055 1.975 371.105 2.025 ;
      RECT 370.935 1.975 370.985 2.025 ;
      RECT 370.815 1.975 370.865 2.025 ;
      RECT 370.695 1.975 370.745 2.025 ;
      RECT 370.575 1.975 370.625 2.025 ;
      RECT 370.455 1.975 370.505 2.025 ;
      RECT 370.335 1.975 370.385 2.025 ;
      RECT 370.215 1.975 370.265 2.025 ;
      RECT 370.095 1.975 370.145 2.025 ;
      RECT 369.975 1.975 370.025 2.025 ;
      RECT 369.855 1.975 369.905 2.025 ;
      RECT 369.735 1.975 369.785 2.025 ;
      RECT 369.615 1.975 369.665 2.025 ;
      RECT 369.495 1.975 369.545 2.025 ;
      RECT 369.375 1.975 369.425 2.025 ;
      RECT 369.255 1.975 369.305 2.025 ;
      RECT 369.135 1.975 369.185 2.025 ;
      RECT 369.015 1.975 369.065 2.025 ;
      RECT 368.895 1.975 368.945 2.025 ;
      RECT 368.775 1.975 368.825 2.025 ;
      RECT 368.655 1.975 368.705 2.025 ;
      RECT 368.535 1.975 368.585 2.025 ;
      RECT 305.415 1.975 305.465 2.025 ;
      RECT 305.295 1.975 305.345 2.025 ;
      RECT 305.175 1.975 305.225 2.025 ;
      RECT 305.055 1.975 305.105 2.025 ;
      RECT 304.935 1.975 304.985 2.025 ;
      RECT 304.815 1.975 304.865 2.025 ;
      RECT 304.695 1.975 304.745 2.025 ;
      RECT 304.575 1.975 304.625 2.025 ;
      RECT 304.455 1.975 304.505 2.025 ;
      RECT 304.335 1.975 304.385 2.025 ;
      RECT 304.215 1.975 304.265 2.025 ;
      RECT 304.095 1.975 304.145 2.025 ;
      RECT 303.975 1.975 304.025 2.025 ;
      RECT 303.855 1.975 303.905 2.025 ;
      RECT 303.735 1.975 303.785 2.025 ;
      RECT 303.615 1.975 303.665 2.025 ;
      RECT 303.495 1.975 303.545 2.025 ;
      RECT 303.375 1.975 303.425 2.025 ;
      RECT 303.255 1.975 303.305 2.025 ;
      RECT 303.135 1.975 303.185 2.025 ;
      RECT 303.015 1.975 303.065 2.025 ;
      RECT 302.895 1.975 302.945 2.025 ;
      RECT 302.775 1.975 302.825 2.025 ;
      RECT 302.655 1.975 302.705 2.025 ;
      RECT 302.535 1.975 302.585 2.025 ;
      RECT 241.415 1.975 241.465 2.025 ;
      RECT 241.295 1.975 241.345 2.025 ;
      RECT 241.175 1.975 241.225 2.025 ;
      RECT 241.055 1.975 241.105 2.025 ;
      RECT 240.935 1.975 240.985 2.025 ;
      RECT 240.815 1.975 240.865 2.025 ;
      RECT 240.695 1.975 240.745 2.025 ;
      RECT 240.575 1.975 240.625 2.025 ;
      RECT 240.455 1.975 240.505 2.025 ;
      RECT 240.335 1.975 240.385 2.025 ;
      RECT 240.215 1.975 240.265 2.025 ;
      RECT 240.095 1.975 240.145 2.025 ;
      RECT 239.975 1.975 240.025 2.025 ;
      RECT 239.855 1.975 239.905 2.025 ;
      RECT 239.735 1.975 239.785 2.025 ;
      RECT 239.615 1.975 239.665 2.025 ;
      RECT 239.495 1.975 239.545 2.025 ;
      RECT 239.375 1.975 239.425 2.025 ;
      RECT 239.255 1.975 239.305 2.025 ;
      RECT 239.135 1.975 239.185 2.025 ;
      RECT 239.015 1.975 239.065 2.025 ;
      RECT 238.895 1.975 238.945 2.025 ;
      RECT 238.775 1.975 238.825 2.025 ;
      RECT 238.655 1.975 238.705 2.025 ;
      RECT 238.535 1.975 238.585 2.025 ;
      RECT 171.415 1.975 171.465 2.025 ;
      RECT 171.295 1.975 171.345 2.025 ;
      RECT 171.175 1.975 171.225 2.025 ;
      RECT 171.055 1.975 171.105 2.025 ;
      RECT 170.935 1.975 170.985 2.025 ;
      RECT 170.815 1.975 170.865 2.025 ;
      RECT 170.695 1.975 170.745 2.025 ;
      RECT 170.575 1.975 170.625 2.025 ;
      RECT 170.455 1.975 170.505 2.025 ;
      RECT 170.335 1.975 170.385 2.025 ;
      RECT 170.215 1.975 170.265 2.025 ;
      RECT 170.095 1.975 170.145 2.025 ;
      RECT 169.975 1.975 170.025 2.025 ;
      RECT 169.855 1.975 169.905 2.025 ;
      RECT 169.735 1.975 169.785 2.025 ;
      RECT 169.615 1.975 169.665 2.025 ;
      RECT 169.495 1.975 169.545 2.025 ;
      RECT 169.375 1.975 169.425 2.025 ;
      RECT 169.255 1.975 169.305 2.025 ;
      RECT 169.135 1.975 169.185 2.025 ;
      RECT 169.015 1.975 169.065 2.025 ;
      RECT 168.895 1.975 168.945 2.025 ;
      RECT 168.775 1.975 168.825 2.025 ;
      RECT 168.655 1.975 168.705 2.025 ;
      RECT 168.535 1.975 168.585 2.025 ;
      RECT 105.415 1.975 105.465 2.025 ;
      RECT 105.295 1.975 105.345 2.025 ;
      RECT 105.175 1.975 105.225 2.025 ;
      RECT 105.055 1.975 105.105 2.025 ;
      RECT 104.935 1.975 104.985 2.025 ;
      RECT 104.815 1.975 104.865 2.025 ;
      RECT 104.695 1.975 104.745 2.025 ;
      RECT 104.575 1.975 104.625 2.025 ;
      RECT 104.455 1.975 104.505 2.025 ;
      RECT 104.335 1.975 104.385 2.025 ;
      RECT 104.215 1.975 104.265 2.025 ;
      RECT 104.095 1.975 104.145 2.025 ;
      RECT 103.975 1.975 104.025 2.025 ;
      RECT 103.855 1.975 103.905 2.025 ;
      RECT 103.735 1.975 103.785 2.025 ;
      RECT 103.615 1.975 103.665 2.025 ;
      RECT 103.495 1.975 103.545 2.025 ;
      RECT 103.375 1.975 103.425 2.025 ;
      RECT 103.255 1.975 103.305 2.025 ;
      RECT 103.135 1.975 103.185 2.025 ;
      RECT 103.015 1.975 103.065 2.025 ;
      RECT 102.895 1.975 102.945 2.025 ;
      RECT 102.775 1.975 102.825 2.025 ;
      RECT 102.655 1.975 102.705 2.025 ;
      RECT 102.535 1.975 102.585 2.025 ;
      RECT 41.415 1.975 41.465 2.025 ;
      RECT 41.295 1.975 41.345 2.025 ;
      RECT 41.175 1.975 41.225 2.025 ;
      RECT 41.055 1.975 41.105 2.025 ;
      RECT 40.935 1.975 40.985 2.025 ;
      RECT 40.815 1.975 40.865 2.025 ;
      RECT 40.695 1.975 40.745 2.025 ;
      RECT 40.575 1.975 40.625 2.025 ;
      RECT 40.455 1.975 40.505 2.025 ;
      RECT 40.335 1.975 40.385 2.025 ;
      RECT 40.215 1.975 40.265 2.025 ;
      RECT 40.095 1.975 40.145 2.025 ;
      RECT 39.975 1.975 40.025 2.025 ;
      RECT 39.855 1.975 39.905 2.025 ;
      RECT 39.735 1.975 39.785 2.025 ;
      RECT 39.615 1.975 39.665 2.025 ;
      RECT 39.495 1.975 39.545 2.025 ;
      RECT 39.375 1.975 39.425 2.025 ;
      RECT 39.255 1.975 39.305 2.025 ;
      RECT 39.135 1.975 39.185 2.025 ;
      RECT 39.015 1.975 39.065 2.025 ;
      RECT 38.895 1.975 38.945 2.025 ;
      RECT 38.775 1.975 38.825 2.025 ;
      RECT 38.655 1.975 38.705 2.025 ;
      RECT 38.535 1.975 38.585 2.025 ;
    LAYER M9 ;
      RECT 0.5 0.5 1638.412 468.316 ;
    LAYER MRDL ;
      RECT 2 2 1636.912 466.816 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 468.816 1638.912 468.816 1638.912 0 ;
  END
END bit_top

END LIBRARY
