class apb_scoreboard extends uvm_scoreboard;

endclass
