`ifndef TR_FILE_LIST__SV 
`define TR_FILE_LIST__SV



`include "btcoin.sv"

 `include "btcoin_seq_sequence_library.sv"
`endif