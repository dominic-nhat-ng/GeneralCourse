class my_sequence extends uvm_sequence #(transaction);

    `uvm_component_object(my_sequence)   
    


endclass
